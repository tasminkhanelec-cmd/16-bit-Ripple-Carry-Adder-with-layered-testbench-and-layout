constraint weight {
    A dist {
      [0    : 63]       :/ A_weights[0],
      [64   : 127]      :/ A_weights[1],
      [128  : 191]      :/ A_weights[2],
      [192  : 255]      :/ A_weights[3],
      [256  : 319]      :/ A_weights[4],
      [320  : 383]      :/ A_weights[5],
      [384  : 447]      :/ A_weights[6],
      [448  : 511]      :/ A_weights[7],
      [512  : 575]      :/ A_weights[8],
      [576  : 639]      :/ A_weights[9],
      [640  : 703]      :/ A_weights[10],
      [704  : 767]      :/ A_weights[11],
      [768  : 831]      :/ A_weights[12],
      [832  : 895]      :/ A_weights[13],
      [896  : 959]      :/ A_weights[14],
      [960  : 1023]     :/ A_weights[15],
      [1024 : 1087]     :/ A_weights[16],
      [1088 : 1151]     :/ A_weights[17],
      [1152 : 1215]     :/ A_weights[18],
      [1216 : 1279]     :/ A_weights[19],
      [1280 : 1343]     :/ A_weights[20],
      [1344 : 1407]     :/ A_weights[21],
      [1408 : 1471]     :/ A_weights[22],
      [1472 : 1535]     :/ A_weights[23],
      [1536 : 1599]     :/ A_weights[24],
      [1600 : 1663]     :/ A_weights[25],
      [1664 : 1727]     :/ A_weights[26],
      [1728 : 1791]     :/ A_weights[27],
      [1792 : 1855]     :/ A_weights[28],
      [1856 : 1919]     :/ A_weights[29],
      [1920 : 1983]     :/ A_weights[30],
      [1984 : 2047]     :/ A_weights[31],
      [2048 : 2111]     :/ A_weights[32],
      [2112 : 2175]     :/ A_weights[33],
      [2176 : 2239]     :/ A_weights[34],
      [2240 : 2303]     :/ A_weights[35],
      [2304 : 2367]     :/ A_weights[36],
      [2368 : 2431]     :/ A_weights[37],
      [2432 : 2495]     :/ A_weights[38],
      [2496 : 2559]     :/ A_weights[39],
      [2560 : 2623]     :/ A_weights[40],
      [2624 : 2687]     :/ A_weights[41],
      [2688 : 2751]     :/ A_weights[42],
      [2752 : 2815]     :/ A_weights[43],
      [2816 : 2879]     :/ A_weights[44],
      [2880 : 2943]     :/ A_weights[45],
      [2944 : 3007]     :/ A_weights[46],
      [3008 : 3071]     :/ A_weights[47],
      [3072 : 3135]     :/ A_weights[48],
      [3136 : 3199]     :/ A_weights[49],
      [3200 : 3263]     :/ A_weights[50],
      [3264 : 3327]     :/ A_weights[51],
      [3328 : 3391]     :/ A_weights[52],
      [3392 : 3455]     :/ A_weights[53],
      [3456 : 3519]     :/ A_weights[54],
      [3520 : 3583]     :/ A_weights[55],
      [3584 : 3647]     :/ A_weights[56],
      [3648 : 3711]     :/ A_weights[57],
      [3712 : 3775]     :/ A_weights[58],
      [3776 : 3839]     :/ A_weights[59],
      [3840 : 3903]     :/ A_weights[60],
      [3904 : 3967]     :/ A_weights[61],
      [3968 : 4031]     :/ A_weights[62],
      [4032 : 4095]     :/ A_weights[63],
      [4096 : 4159]     :/ A_weights[64],
      [4160 : 4223]     :/ A_weights[65],
      [4224 : 4287]     :/ A_weights[66],
      [4288 : 4351]     :/ A_weights[67],
      [4352 : 4415]     :/ A_weights[68],
      [4416 : 4479]     :/ A_weights[69],
      [4480 : 4543]     :/ A_weights[70],
      [4544 : 4607]     :/ A_weights[71],
      [4608 : 4671]     :/ A_weights[72],
      [4672 : 4735]     :/ A_weights[73],
      [4736 : 4799]     :/ A_weights[74],
      [4800 : 4863]     :/ A_weights[75],
      [4864 : 4927]     :/ A_weights[76],
      [4928 : 4991]     :/ A_weights[77],
      [4992 : 5055]     :/ A_weights[78],
      [5056 : 5119]     :/ A_weights[79],
      [5120 : 5183]     :/ A_weights[80],
      [5184 : 5247]     :/ A_weights[81],
      [5248 : 5311]     :/ A_weights[82],
      [5312 : 5375]     :/ A_weights[83],
      [5376 : 5439]     :/ A_weights[84],
      [5440 : 5503]     :/ A_weights[85],
      [5504 : 5567]     :/ A_weights[86],
      [5568 : 5631]     :/ A_weights[87],
      [5632 : 5695]     :/ A_weights[88],
      [5696 : 5759]     :/ A_weights[89],
      [5760 : 5823]     :/ A_weights[90],
      [5824 : 5887]     :/ A_weights[91],
      [5888 : 5951]     :/ A_weights[92],
      [5952 : 6015]     :/ A_weights[93],
      [6016 : 6079]     :/ A_weights[94],
      [6080 : 6143]     :/ A_weights[95],
      [6144 : 6207]     :/ A_weights[96],
      [6208 : 6271]     :/ A_weights[97],
      [6272 : 6335]     :/ A_weights[98],
      [6336 : 6399]     :/ A_weights[99],
      [6400 : 6463]     :/ A_weights[100],
      [6464 : 6527]     :/ A_weights[101],
      [6528 : 6591]     :/ A_weights[102],
      [6592 : 6655]     :/ A_weights[103],
      [6656 : 6719]     :/ A_weights[104],
      [6720 : 6783]     :/ A_weights[105],
      [6784 : 6847]     :/ A_weights[106],
      [6848 : 6911]     :/ A_weights[107],
      [6912 : 6975]     :/ A_weights[108],
      [6976 : 7039]     :/ A_weights[109],
      [7040 : 7103]     :/ A_weights[110],
      [7104 : 7167]     :/ A_weights[111],
      [7168 : 7231]     :/ A_weights[112],
      [7232 : 7295]     :/ A_weights[113],
      [7296 : 7359]     :/ A_weights[114],
      [7360 : 7423]     :/ A_weights[115],
      [7424 : 7487]     :/ A_weights[116],
      [7488 : 7551]     :/ A_weights[117],
      [7552 : 7615]     :/ A_weights[118],
      [7616 : 7679]     :/ A_weights[119],
      [7680 : 7743]     :/ A_weights[120],
      [7744 : 7807]     :/ A_weights[121],
      [7808 : 7871]     :/ A_weights[122],
      [7872 : 7935]     :/ A_weights[123],
      [7936 : 7999]     :/ A_weights[124],
      [8000 : 8063]     :/ A_weights[125],
      [8064 : 8127]     :/ A_weights[126],
      [8128 : 8191]     :/ A_weights[127],
      [8192 : 8255]     :/ A_weights[128],
      [8256 : 8319]     :/ A_weights[129],
      [8320 : 8383]     :/ A_weights[130],
      [8384 : 8447]     :/ A_weights[131],
      [8448 : 8511]     :/ A_weights[132],
      [8512 : 8575]     :/ A_weights[133],
      [8576 : 8639]     :/ A_weights[134],
      [8640 : 8703]     :/ A_weights[135],
      [8704 : 8767]     :/ A_weights[136],
      [8768 : 8831]     :/ A_weights[137],
      [8832 : 8895]     :/ A_weights[138],
      [8896 : 8959]     :/ A_weights[139],
      [8960 : 9023]     :/ A_weights[140],
      [9024 : 9087]     :/ A_weights[141],
      [9088 : 9151]     :/ A_weights[142],
      [9152 : 9215]     :/ A_weights[143],
      [9216 : 9279]     :/ A_weights[144],
      [9280 : 9343]     :/ A_weights[145],
      [9344 : 9407]     :/ A_weights[146],
      [9408 : 9471]     :/ A_weights[147],
      [9472 : 9535]     :/ A_weights[148],
      [9536 : 9599]     :/ A_weights[149],
      [9600 : 9663]     :/ A_weights[150],
      [9664 : 9727]     :/ A_weights[151],
      [9728 : 9791]     :/ A_weights[152],
      [9792 : 9855]     :/ A_weights[153],
      [9856 : 9919]     :/ A_weights[154],
      [9920 : 9983]     :/ A_weights[155],
      [9984 : 10047]    :/ A_weights[156],
      [10048 : 10111]   :/ A_weights[157],
      [10112 : 10175]   :/ A_weights[158],
      [10176 : 10239]   :/ A_weights[159],
      [10240 : 10303]   :/ A_weights[160],
      [10304 : 10367]   :/ A_weights[161],
      [10368 : 10431]   :/ A_weights[162],
      [10432 : 10495]   :/ A_weights[163],
      [10496 : 10559]   :/ A_weights[164],
      [10560 : 10623]   :/ A_weights[165],
      [10624 : 10687]   :/ A_weights[166],
      [10688 : 10751]   :/ A_weights[167],
      [10752 : 10815]   :/ A_weights[168],
      [10816 : 10879]   :/ A_weights[169],
      [10880 : 10943]   :/ A_weights[170],
      [10944 : 11007]   :/ A_weights[171],
      [11008 : 11071]   :/ A_weights[172],
      [11072 : 11135]   :/ A_weights[173],
      [11136 : 11199]   :/ A_weights[174],
      [11200 : 11263]   :/ A_weights[175],
      [11264 : 11327]   :/ A_weights[176],
      [11328 : 11391]   :/ A_weights[177],
      [11392 : 11455]   :/ A_weights[178],
      [11456 : 11519]   :/ A_weights[179],
      [11520 : 11583]   :/ A_weights[180],
      [11584 : 11647]   :/ A_weights[181],
      [11648 : 11711]   :/ A_weights[182],
      [11712 : 11775]   :/ A_weights[183],
      [11776 : 11839]   :/ A_weights[184],
      [11840 : 11903]   :/ A_weights[185],
      [11904 : 11967]   :/ A_weights[186],
      [11968 : 12031]   :/ A_weights[187],
      [12032 : 12095]   :/ A_weights[188],
      [12096 : 12159]   :/ A_weights[189],
      [12160 : 12223]   :/ A_weights[190],
      [12224 : 12287]   :/ A_weights[191],
      [12288 : 12351]   :/ A_weights[192],
      [12352 : 12415]   :/ A_weights[193],
      [12416 : 12479]   :/ A_weights[194],
      [12480 : 12543]   :/ A_weights[195],
      [12544 : 12607]   :/ A_weights[196],
      [12608 : 12671]   :/ A_weights[197],
      [12672 : 12735]   :/ A_weights[198],
      [12736 : 12799]   :/ A_weights[199],
      [12800 : 12863]   :/ A_weights[200],
      [12864 : 12927]   :/ A_weights[201],
      [12928 : 12991]   :/ A_weights[202],
      [12992 : 13055]   :/ A_weights[203],
      [13056 : 13119]   :/ A_weights[204],
      [13120 : 13183]   :/ A_weights[205],
      [13184 : 13247]   :/ A_weights[206],
      [13248 : 13311]   :/ A_weights[207],
      [13312 : 13375]   :/ A_weights[208],
      [13376 : 13439]   :/ A_weights[209],
      [13440 : 13503]   :/ A_weights[210],
      [13504 : 13567]   :/ A_weights[211],
      [13568 : 13631]   :/ A_weights[212],
      [13632 : 13695]   :/ A_weights[213],
      [13696 : 13759]   :/ A_weights[214],
      [13760 : 13823]   :/ A_weights[215],
      [13824 : 13887]   :/ A_weights[216],
      [13888 : 13951]   :/ A_weights[217],
      [13952 : 14015]   :/ A_weights[218],
      [14016 : 14079]   :/ A_weights[219],
      [14080 : 14143]   :/ A_weights[220],
      [14144 : 14207]   :/ A_weights[221],
      [14208 : 14271]   :/ A_weights[222],
      [14272 : 14335]   :/ A_weights[223],
      [14336 : 14399]   :/ A_weights[224],
      [14400 : 14463]   :/ A_weights[225],
      [14464 : 14527]   :/ A_weights[226],
      [14528 : 14591]   :/ A_weights[227],
      [14592 : 14655]   :/ A_weights[228],
      [14656 : 14719]   :/ A_weights[229],
      [14720 : 14783]   :/ A_weights[230],
      [14784 : 14847]   :/ A_weights[231],
      [14848 : 14911]   :/ A_weights[232],
      [14912 : 14975]   :/ A_weights[233],
      [14976 : 15039]   :/ A_weights[234],
      [15040 : 15103]   :/ A_weights[235],
      [15104 : 15167]   :/ A_weights[236],
      [15168 : 15231]   :/ A_weights[237],
      [15232 : 15295]   :/ A_weights[238],
      [15296 : 15359]   :/ A_weights[239],
      [15360 : 15423]   :/ A_weights[240],
      [15424 : 15487]   :/ A_weights[241],
      [15488 : 15551]   :/ A_weights[242],
      [15552 : 15615]   :/ A_weights[243],
      [15616 : 15679]   :/ A_weights[244],
      [15680 : 15743]   :/ A_weights[245],
      [15744 : 15807]   :/ A_weights[246],
      [15808 : 15871]   :/ A_weights[247],
      [15872 : 15935]   :/ A_weights[248],
      [15936 : 15999]   :/ A_weights[249],
      [16000 : 16063]   :/ A_weights[250],
      [16064 : 16127]   :/ A_weights[251],
      [16128 : 16191]   :/ A_weights[252],
      [16192 : 16255]   :/ A_weights[253],
      [16256 : 16319]   :/ A_weights[254],
      [16320 : 16383]   :/ A_weights[255],
      [16384 : 16447]   :/ A_weights[256],
      [16448 : 16511]   :/ A_weights[257],
      [16512 : 16575]   :/ A_weights[258],
      [16576 : 16639]   :/ A_weights[259],
      [16640 : 16703]   :/ A_weights[260],
      [16704 : 16767]   :/ A_weights[261],
      [16768 : 16831]   :/ A_weights[262],
      [16832 : 16895]   :/ A_weights[263],
      [16896 : 16959]   :/ A_weights[264],
      [16960 : 17023]   :/ A_weights[265],
      [17024 : 17087]   :/ A_weights[266],
      [17088 : 17151]   :/ A_weights[267],
      [17152 : 17215]   :/ A_weights[268],
      [17216 : 17279]   :/ A_weights[269],
      [17280 : 17343]   :/ A_weights[270],
      [17344 : 17407]   :/ A_weights[271],
      [17408 : 17471]   :/ A_weights[272],
      [17472 : 17535]   :/ A_weights[273],
      [17536 : 17599]   :/ A_weights[274],
      [17600 : 17663]   :/ A_weights[275],
      [17664 : 17727]   :/ A_weights[276],
      [17728 : 17791]   :/ A_weights[277],
      [17792 : 17855]   :/ A_weights[278],
      [17856 : 17919]   :/ A_weights[279],
      [17920 : 17983]   :/ A_weights[280],
      [17984 : 18047]   :/ A_weights[281],
      [18048 : 18111]   :/ A_weights[282],
      [18112 : 18175]   :/ A_weights[283],
      [18176 : 18239]   :/ A_weights[284],
      [18240 : 18303]   :/ A_weights[285],
      [18304 : 18367]   :/ A_weights[286],
      [18368 : 18431]   :/ A_weights[287],
      [18432 : 18495]   :/ A_weights[288],
      [18496 : 18559]   :/ A_weights[289],
      [18560 : 18623]   :/ A_weights[290],
      [18624 : 18687]   :/ A_weights[291],
      [18688 : 18751]   :/ A_weights[292],
      [18752 : 18815]   :/ A_weights[293],
      [18816 : 18879]   :/ A_weights[294],
      [18880 : 18943]   :/ A_weights[295],
      [18944 : 19007]   :/ A_weights[296],
      [19008 : 19071]   :/ A_weights[297],
      [19072 : 19135]   :/ A_weights[298],
      [19136 : 19199]   :/ A_weights[299],
      [19200 : 19263]   :/ A_weights[300],
      [19264 : 19327]   :/ A_weights[301],
      [19328 : 19391]   :/ A_weights[302],
      [19392 : 19455]   :/ A_weights[303],
      [19456 : 19519]   :/ A_weights[304],
      [19520 : 19583]   :/ A_weights[305],
      [19584 : 19647]   :/ A_weights[306],
      [19648 : 19711]   :/ A_weights[307],
      [19712 : 19775]   :/ A_weights[308],
      [19776 : 19839]   :/ A_weights[309],
      [19840 : 19903]   :/ A_weights[310],
      [19904 : 19967]   :/ A_weights[311],
      [19968 : 20031]   :/ A_weights[312],
      [20032 : 20095]   :/ A_weights[313],
      [20096 : 20159]   :/ A_weights[314],
      [20160 : 20223]   :/ A_weights[315],
      [20224 : 20287]   :/ A_weights[316],
      [20288 : 20351]   :/ A_weights[317],
      [20352 : 20415]   :/ A_weights[318],
      [20416 : 20479]   :/ A_weights[319],
      [20480 : 20543]   :/ A_weights[320],
      [20544 : 20607]   :/ A_weights[321],
      [20608 : 20671]   :/ A_weights[322],
      [20672 : 20735]   :/ A_weights[323],
      [20736 : 20799]   :/ A_weights[324],
      [20800 : 20863]   :/ A_weights[325],
      [20864 : 20927]   :/ A_weights[326],
      [20928 : 20991]   :/ A_weights[327],
      [20992 : 21055]   :/ A_weights[328],
      [21056 : 21119]   :/ A_weights[329],
      [21120 : 21183]   :/ A_weights[330],
      [21184 : 21247]   :/ A_weights[331],
      [21248 : 21311]   :/ A_weights[332],
      [21312 : 21375]   :/ A_weights[333],
      [21376 : 21439]   :/ A_weights[334],
      [21440 : 21503]   :/ A_weights[335],
      [21504 : 21567]   :/ A_weights[336],
      [21568 : 21631]   :/ A_weights[337],
      [21632 : 21695]   :/ A_weights[338],
      [21696 : 21759]   :/ A_weights[339],
      [21760 : 21823]   :/ A_weights[340],
      [21824 : 21887]   :/ A_weights[341],
      [21888 : 21951]   :/ A_weights[342],
      [21952 : 22015]   :/ A_weights[343],
      [22016 : 22079]   :/ A_weights[344],
      [22080 : 22143]   :/ A_weights[345],
      [22144 : 22207]   :/ A_weights[346],
      [22208 : 22271]   :/ A_weights[347],
      [22272 : 22335]   :/ A_weights[348],
      [22336 : 22399]   :/ A_weights[349],
      [22400 : 22463]   :/ A_weights[350],
      [22464 : 22527]   :/ A_weights[351],
      [22528 : 22591]   :/ A_weights[352],
      [22592 : 22655]   :/ A_weights[353],
      [22656 : 22719]   :/ A_weights[354],
      [22720 : 22783]   :/ A_weights[355],
      [22784 : 22847]   :/ A_weights[356],
      [22848 : 22911]   :/ A_weights[357],
      [22912 : 22975]   :/ A_weights[358],
      [22976 : 23039]   :/ A_weights[359],
      [23040 : 23103]   :/ A_weights[360],
      [23104 : 23167]   :/ A_weights[361],
      [23168 : 23231]   :/ A_weights[362],
      [23232 : 23295]   :/ A_weights[363],
      [23296 : 23359]   :/ A_weights[364],
      [23360 : 23423]   :/ A_weights[365],
      [23424 : 23487]   :/ A_weights[366],
      [23488 : 23551]   :/ A_weights[367],
      [23552 : 23615]   :/ A_weights[368],
      [23616 : 23679]   :/ A_weights[369],
      [23680 : 23743]   :/ A_weights[370],
      [23744 : 23807]   :/ A_weights[371],
      [23808 : 23871]   :/ A_weights[372],
      [23872 : 23935]   :/ A_weights[373],
      [23936 : 23999]   :/ A_weights[374],
      [24000 : 24063]   :/ A_weights[375],
      [24064 : 24127]   :/ A_weights[376],
      [24128 : 24191]   :/ A_weights[377],
      [24192 : 24255]   :/ A_weights[378],
      [24256 : 24319]   :/ A_weights[379],
      [24320 : 24383]   :/ A_weights[380],
      [24384 : 24447]   :/ A_weights[381],
      [24448 : 24511]   :/ A_weights[382],
      [24512 : 24575]   :/ A_weights[383],
      [24576 : 24639]   :/ A_weights[384],
      [24640 : 24703]   :/ A_weights[385],
      [24704 : 24767]   :/ A_weights[386],
      [24768 : 24831]   :/ A_weights[387],
      [24832 : 24895]   :/ A_weights[388],
      [24896 : 24959]   :/ A_weights[389],
      [24960 : 25023]   :/ A_weights[390],
      [25024 : 25087]   :/ A_weights[391],
      [25088 : 25151]   :/ A_weights[392],
      [25152 : 25215]   :/ A_weights[393],
      [25216 : 25279]   :/ A_weights[394],
      [25280 : 25343]   :/ A_weights[395],
      [25344 : 25407]   :/ A_weights[396],
      [25408 : 25471]   :/ A_weights[397],
      [25472 : 25535]   :/ A_weights[398],
      [25536 : 25599]   :/ A_weights[399],
      [25600 : 25663]   :/ A_weights[400],
      [25664 : 25727]   :/ A_weights[401],
      [25728 : 25791]   :/ A_weights[402],
      [25792 : 25855]   :/ A_weights[403],
      [25856 : 25919]   :/ A_weights[404],
      [25920 : 25983]   :/ A_weights[405],
      [25984 : 26047]   :/ A_weights[406],
      [26048 : 26111]   :/ A_weights[407],
      [26112 : 26175]   :/ A_weights[408],
      [26176 : 26239]   :/ A_weights[409],
      [26240 : 26303]   :/ A_weights[410],
      [26304 : 26367]   :/ A_weights[411],
      [26368 : 26431]   :/ A_weights[412],
      [26432 : 26495]   :/ A_weights[413],
      [26496 : 26559]   :/ A_weights[414],
      [26560 : 26623]   :/ A_weights[415],
      [26624 : 26687]   :/ A_weights[416],
      [26688 : 26751]   :/ A_weights[417],
      [26752 : 26815]   :/ A_weights[418],
      [26816 : 26879]   :/ A_weights[419],
      [26880 : 26943]   :/ A_weights[420],
      [26944 : 27007]   :/ A_weights[421],
      [27008 : 27071]   :/ A_weights[422],
      [27072 : 27135]   :/ A_weights[423],
      [27136 : 27199]   :/ A_weights[424],
      [27200 : 27263]   :/ A_weights[425],
      [27264 : 27327]   :/ A_weights[426],
      [27328 : 27391]   :/ A_weights[427],
      [27392 : 27455]   :/ A_weights[428],
      [27456 : 27519]   :/ A_weights[429],
      [27520 : 27583]   :/ A_weights[430],
      [27584 : 27647]   :/ A_weights[431],
      [27648 : 27711]   :/ A_weights[432],
      [27712 : 27775]   :/ A_weights[433],
      [27776 : 27839]   :/ A_weights[434],
      [27840 : 27903]   :/ A_weights[435],
      [27904 : 27967]   :/ A_weights[436],
      [27968 : 28031]   :/ A_weights[437],
      [28032 : 28095]   :/ A_weights[438],
      [28096 : 28159]   :/ A_weights[439],
      [28160 : 28223]   :/ A_weights[440],
      [28224 : 28287]   :/ A_weights[441],
      [28288 : 28351]   :/ A_weights[442],
      [28352 : 28415]   :/ A_weights[443],
      [28416 : 28479]   :/ A_weights[444],
      [28480 : 28543]   :/ A_weights[445],
      [28544 : 28607]   :/ A_weights[446],
      [28608 : 28671]   :/ A_weights[447],
      [28672 : 28735]   :/ A_weights[448],
      [28736 : 28799]   :/ A_weights[449],
      [28800 : 28863]   :/ A_weights[450],
      [28864 : 28927]   :/ A_weights[451],
      [28928 : 28991]   :/ A_weights[452],
      [28992 : 29055]   :/ A_weights[453],
      [29056 : 29119]   :/ A_weights[454],
      [29120 : 29183]   :/ A_weights[455],
      [29184 : 29247]   :/ A_weights[456],
      [29248 : 29311]   :/ A_weights[457],
      [29312 : 29375]   :/ A_weights[458],
      [29376 : 29439]   :/ A_weights[459],
      [29440 : 29503]   :/ A_weights[460],
      [29504 : 29567]   :/ A_weights[461],
      [29568 : 29631]   :/ A_weights[462],
      [29632 : 29695]   :/ A_weights[463],
      [29696 : 29759]   :/ A_weights[464],
      [29760 : 29823]   :/ A_weights[465],
      [29824 : 29887]   :/ A_weights[466],
      [29888 : 29951]   :/ A_weights[467],
      [29952 : 30015]   :/ A_weights[468],
      [30016 : 30079]   :/ A_weights[469],
      [30080 : 30143]   :/ A_weights[470],
      [30144 : 30207]   :/ A_weights[471],
      [30208 : 30271]   :/ A_weights[472],
      [30272 : 30335]   :/ A_weights[473],
      [30336 : 30399]   :/ A_weights[474],
      [30400 : 30463]   :/ A_weights[475],
      [30464 : 30527]   :/ A_weights[476],
      [30528 : 30591]   :/ A_weights[477],
      [30592 : 30655]   :/ A_weights[478],
      [30656 : 30719]   :/ A_weights[479],
      [30720 : 30783]   :/ A_weights[480],
      [30784 : 30847]   :/ A_weights[481],
      [30848 : 30911]   :/ A_weights[482],
      [30912 : 30975]   :/ A_weights[483],
      [30976 : 31039]   :/ A_weights[484],
      [31040 : 31103]   :/ A_weights[485],
      [31104 : 31167]   :/ A_weights[486],
      [31168 : 31231]   :/ A_weights[487],
      [31232 : 31295]   :/ A_weights[488],
      [31296 : 31359]   :/ A_weights[489],
      [31360 : 31423]   :/ A_weights[490],
      [31424 : 31487]   :/ A_weights[491],
      [31488 : 31551]   :/ A_weights[492],
      [31552 : 31615]   :/ A_weights[493],
      [31616 : 31679]   :/ A_weights[494],
      [31680 : 31743]   :/ A_weights[495],
      [31744 : 31807]   :/ A_weights[496],
      [31808 : 31871]   :/ A_weights[497],
      [31872 : 31935]   :/ A_weights[498],
      [31936 : 31999]   :/ A_weights[499],
      [32000 : 32063]   :/ A_weights[500],      
      [32064 : 32127]   :/ A_weights[501],
      [32128 : 32191]   :/ A_weights[502],
      [32192 : 32255]   :/ A_weights[503],
      [32256 : 32319]   :/ A_weights[504],
      [32320 : 32383]   :/ A_weights[505],
      [32384 : 32447]   :/ A_weights[506],
      [32448 : 32511]   :/ A_weights[507],
      [32512 : 32575]   :/ A_weights[508],
      [32576 : 32639]   :/ A_weights[509],
      [32640 : 32703]   :/ A_weights[510],
      [32704 : 32767]   :/ A_weights[511],
      [32768 : 32831]   :/ A_weights[512],
      [32832 : 32895]   :/ A_weights[513],
      [32896 : 32959]   :/ A_weights[514],
      [32960 : 33023]   :/ A_weights[515],
      [33024 : 33087]   :/ A_weights[516],
      [33088 : 33151]   :/ A_weights[517],
      [33152 : 33215]   :/ A_weights[518],
      [33216 : 33279]   :/ A_weights[519],
      [33280 : 33343]   :/ A_weights[520],
      [33344 : 33407]   :/ A_weights[521],
      [33408 : 33471]   :/ A_weights[522],
      [33472 : 33535]   :/ A_weights[523],
      [33536 : 33599]   :/ A_weights[524],
      [33600 : 33663]   :/ A_weights[525],
      [33664 : 33727]   :/ A_weights[526],
      [33728 : 33791]   :/ A_weights[527],
      [33792 : 33855]   :/ A_weights[528],
      [33856 : 33919]   :/ A_weights[529],
      [33920 : 33983]   :/ A_weights[530],
      [33984 : 34047]   :/ A_weights[531],
      [34048 : 34111]   :/ A_weights[532],
      [34112 : 34175]   :/ A_weights[533],
      [34176 : 34239]   :/ A_weights[534],
      [34240 : 34303]   :/ A_weights[535],
      [34304 : 34367]   :/ A_weights[536],
      [34368 : 34431]   :/ A_weights[537],
      [34432 : 34495]   :/ A_weights[538],
      [34496 : 34559]   :/ A_weights[539],
      [34560 : 34623]   :/ A_weights[540],
      [34624 : 34687]   :/ A_weights[541],
      [34688 : 34751]   :/ A_weights[542],
      [34752 : 34815]   :/ A_weights[543],
      [34816 : 34879]   :/ A_weights[544],
      [34880 : 34943]   :/ A_weights[545],
      [34944 : 35007]   :/ A_weights[546],
      [35008 : 35071]   :/ A_weights[547],
      [35072 : 35135]   :/ A_weights[548],
      [35136 : 35199]   :/ A_weights[549],
      [35200 : 35263]   :/ A_weights[550],
      [35264 : 35327]   :/ A_weights[551],
      [35328 : 35391]   :/ A_weights[552],
      [35392 : 35455]   :/ A_weights[553],
      [35456 : 35519]   :/ A_weights[554],
      [35520 : 35583]   :/ A_weights[555],
      [35584 : 35647]   :/ A_weights[556],
      [35648 : 35711]   :/ A_weights[557],
      [35712 : 35775]   :/ A_weights[558],
      [35776 : 35839]   :/ A_weights[559],
      [35840 : 35903]   :/ A_weights[560],
      [35904 : 35967]   :/ A_weights[561],
      [35968 : 36031]   :/ A_weights[562],
      [36032 : 36095]   :/ A_weights[563],
      [36096 : 36159]   :/ A_weights[564],
      [36160 : 36223]   :/ A_weights[565],
      [36224 : 36287]   :/ A_weights[566],
      [36288 : 36351]   :/ A_weights[567],
      [36352 : 36415]   :/ A_weights[568],
      [36416 : 36479]   :/ A_weights[569],
      [36480 : 36543]   :/ A_weights[570],
      [36544 : 36607]   :/ A_weights[571],
      [36608 : 36671]   :/ A_weights[572],
      [36672 : 36735]   :/ A_weights[573],
      [36736 : 36799]   :/ A_weights[574],
      [36800 : 36863]   :/ A_weights[575],
      [36864 : 36927]   :/ A_weights[576],
      [36928 : 36991]   :/ A_weights[577],
      [36992 : 37055]   :/ A_weights[578],
      [37056 : 37119]   :/ A_weights[579],
      [37120 : 37183]   :/ A_weights[580],
      [37184 : 37247]   :/ A_weights[581],
      [37248 : 37311]   :/ A_weights[582],
      [37312 : 37375]   :/ A_weights[583],
      [37376 : 37439]   :/ A_weights[584],
      [37440 : 37503]   :/ A_weights[585],
      [37504 : 37567]   :/ A_weights[586],
      [37568 : 37631]   :/ A_weights[587],
      [37632 : 37695]   :/ A_weights[588],
      [37696 : 37759]   :/ A_weights[589],
      [37760 : 37823]   :/ A_weights[590],
      [37824 : 37887]   :/ A_weights[591],
      [37888 : 37951]   :/ A_weights[592],
      [37952 : 38015]   :/ A_weights[593],
      [38016 : 38079]   :/ A_weights[594],
      [38080 : 38143]   :/ A_weights[595],
      [38144 : 38207]   :/ A_weights[596],
      [38208 : 38271]   :/ A_weights[597],
      [38272 : 38335]   :/ A_weights[598],
      [38336 : 38399]   :/ A_weights[599],
      [38400 : 38463]   :/ A_weights[600],
      [38464 : 38527]   :/ A_weights[601],
      [38528 : 38591]   :/ A_weights[602],
      [38592 : 38655]   :/ A_weights[603],
      [38656 : 38719]   :/ A_weights[604],
      [38720 : 38783]   :/ A_weights[605],
      [38784 : 38847]   :/ A_weights[606],
      [38848 : 38911]   :/ A_weights[607],
      [38912 : 38975]   :/ A_weights[608],
      [38976 : 39039]   :/ A_weights[609],
      [39040 : 39103]   :/ A_weights[610],
      [39104 : 39167]   :/ A_weights[611],
      [39168 : 39231]   :/ A_weights[612],
      [39232 : 39295]   :/ A_weights[613],
      [39296 : 39359]   :/ A_weights[614],
      [39360 : 39423]   :/ A_weights[615],
      [39424 : 39487]   :/ A_weights[616],
      [39488 : 39551]   :/ A_weights[617],
      [39552 : 39615]   :/ A_weights[618],
      [39616 : 39679]   :/ A_weights[619],
      [39680 : 39743]   :/ A_weights[620],
      [39744 : 39807]   :/ A_weights[621],
      [39808 : 39871]   :/ A_weights[622],
      [39872 : 39935]   :/ A_weights[623],
      [39936 : 39999]   :/ A_weights[624],
      [40000 : 40063]   :/ A_weights[625],
      [40064 : 40127]   :/ A_weights[626],
      [40128 : 40191]   :/ A_weights[627],
      [40192 : 40255]   :/ A_weights[628],
      [40256 : 40319]   :/ A_weights[629],
      [40320 : 40383]   :/ A_weights[630],
      [40384 : 40447]   :/ A_weights[631],
      [40448 : 40511]   :/ A_weights[632],
      [40512 : 40575]   :/ A_weights[633],
      [40576 : 40639]   :/ A_weights[634],
      [40640 : 40703]   :/ A_weights[635],
      [40704 : 40767]   :/ A_weights[636],
      [40768 : 40831]   :/ A_weights[637],
      [40832 : 40895]   :/ A_weights[638],
      [40896 : 40959]   :/ A_weights[639],
      [40960 : 41023]   :/ A_weights[640],
      [41024 : 41087]   :/ A_weights[641],
      [41088 : 41151]   :/ A_weights[642],
      [41152 : 41215]   :/ A_weights[643],
      [41216 : 41279]   :/ A_weights[644],
      [41280 : 41343]   :/ A_weights[645],
      [41344 : 41407]   :/ A_weights[646],
      [41408 : 41471]   :/ A_weights[647],
      [41472 : 41535]   :/ A_weights[648],
      [41536 : 41599]   :/ A_weights[649],
      [41600 : 41663]   :/ A_weights[650],
      [41664 : 41727]   :/ A_weights[651],
      [41728 : 41791]   :/ A_weights[652],
      [41792 : 41855]   :/ A_weights[653],
      [41856 : 41919]   :/ A_weights[654],
      [41920 : 41983]   :/ A_weights[655],
      [41984 : 42047]   :/ A_weights[656],
      [42048 : 42111]   :/ A_weights[657],
      [42112 : 42175]   :/ A_weights[658],
      [42176 : 42239]   :/ A_weights[659],
      [42240 : 42303]   :/ A_weights[660],
      [42304 : 42367]   :/ A_weights[661],
      [42368 : 42431]   :/ A_weights[662],
      [42432 : 42495]   :/ A_weights[663],
      [42496 : 42559]   :/ A_weights[664],
      [42560 : 42623]   :/ A_weights[665],
      [42624 : 42687]   :/ A_weights[666],
      [42688 : 42751]   :/ A_weights[667],
      [42752 : 42815]   :/ A_weights[668],
      [42816 : 42879]   :/ A_weights[669],
      [42880 : 42943]   :/ A_weights[670],
      [42944 : 43007]   :/ A_weights[671],
      [43008 : 43071]   :/ A_weights[672],
      [43072 : 43135]   :/ A_weights[673],
      [43136 : 43199]   :/ A_weights[674],
      [43200 : 43263]   :/ A_weights[675],
      [43264 : 43327]   :/ A_weights[676],
      [43328 : 43391]   :/ A_weights[677],
      [43392 : 43455]   :/ A_weights[678],
      [43456 : 43519]   :/ A_weights[679],
      [43520 : 43583]   :/ A_weights[680],
      [43584 : 43647]   :/ A_weights[681],
      [43648 : 43711]   :/ A_weights[682],
      [43712 : 43775]   :/ A_weights[683],
      [43776 : 43839]   :/ A_weights[684],
      [43840 : 43903]   :/ A_weights[685],
      [43904 : 43967]   :/ A_weights[686],
      [43968 : 44031]   :/ A_weights[687],
      [44032 : 44095]   :/ A_weights[688],
      [44096 : 44159]   :/ A_weights[689],
      [44160 : 44223]   :/ A_weights[690],
      [44224 : 44287]   :/ A_weights[691],
      [44288 : 44351]   :/ A_weights[692],
      [44352 : 44415]   :/ A_weights[693],
      [44416 : 44479]   :/ A_weights[694],
      [44480 : 44543]   :/ A_weights[695],
      [44544 : 44607]   :/ A_weights[696],
      [44608 : 44671]   :/ A_weights[697],
      [44672 : 44735]   :/ A_weights[698],
      [44736 : 44799]   :/ A_weights[699],
      [44800 : 44863]   :/ A_weights[700],
      [44864 : 44927]   :/ A_weights[701],
      [44928 : 44991]   :/ A_weights[702],
      [44992 : 45055]   :/ A_weights[703],
      [45056 : 45119]   :/ A_weights[704],
      [45120 : 45183]   :/ A_weights[705],
      [45184 : 45247]   :/ A_weights[706],
      [45248 : 45311]   :/ A_weights[707],
      [45312 : 45375]   :/ A_weights[708],
      [45376 : 45439]   :/ A_weights[709],
      [45440 : 45503]   :/ A_weights[710],
      [45504 : 45567]   :/ A_weights[711],
      [45568 : 45631]   :/ A_weights[712],
      [45632 : 45695]   :/ A_weights[713],
      [45696 : 45759]   :/ A_weights[714],
      [45760 : 45823]   :/ A_weights[715],
      [45824 : 45887]   :/ A_weights[716],
      [45888 : 45951]   :/ A_weights[717],
      [45952 : 46015]   :/ A_weights[718],
      [46016 : 46079]   :/ A_weights[719],
      [46080 : 46143]   :/ A_weights[720],
      [46144 : 46207]   :/ A_weights[721],
      [46208 : 46271]   :/ A_weights[722],
      [46272 : 46335]   :/ A_weights[723],
      [46336 : 46399]   :/ A_weights[724],
      [46400 : 46463]   :/ A_weights[725],
      [46464 : 46527]   :/ A_weights[726],
      [46528 : 46591]   :/ A_weights[727],
      [46592 : 46655]   :/ A_weights[728],
      [46656 : 46719]   :/ A_weights[729],
      [46720 : 46783]   :/ A_weights[730],
      [46784 : 46847]   :/ A_weights[731],
      [46848 : 46911]   :/ A_weights[732],
      [46912 : 46975]   :/ A_weights[733],
      [46976 : 47039]   :/ A_weights[734],
      [47040 : 47103]   :/ A_weights[735],
      [47104 : 47167]   :/ A_weights[736],
      [47168 : 47231]   :/ A_weights[737],
      [47232 : 47295]   :/ A_weights[738],
      [47296 : 47359]   :/ A_weights[739],
      [47360 : 47423]   :/ A_weights[740],
      [47424 : 47487]   :/ A_weights[741],
      [47488 : 47551]   :/ A_weights[742],
      [47552 : 47615]   :/ A_weights[743],
      [47616 : 47679]   :/ A_weights[744],
      [47680 : 47743]   :/ A_weights[745],
      [47744 : 47807]   :/ A_weights[746],
      [47808 : 47871]   :/ A_weights[747],
      [47872 : 47935]   :/ A_weights[748],
      [47936 : 47999]   :/ A_weights[749],
      [48000 : 48063]   :/ A_weights[750],
      [48064 : 48127]   :/ A_weights[751],
      [48128 : 48191]   :/ A_weights[752],
      [48192 : 48255]   :/ A_weights[753],
      [48256 : 48319]   :/ A_weights[754],
      [48320 : 48383]   :/ A_weights[755],
      [48384 : 48447]   :/ A_weights[756],
      [48448 : 48511]   :/ A_weights[757],
      [48512 : 48575]   :/ A_weights[758],
      [48576 : 48639]   :/ A_weights[759],
      [48640 : 48703]   :/ A_weights[760],
      [48704 : 48767]   :/ A_weights[761],
      [48768 : 48831]   :/ A_weights[762],
      [48832 : 48895]   :/ A_weights[763],
      [48896 : 48959]   :/ A_weights[764],
      [48960 : 49023]   :/ A_weights[765],
      [49024 : 49087]   :/ A_weights[766],
      [49088 : 49151]   :/ A_weights[767],
      [49152 : 49215]   :/ A_weights[768],
      [49216 : 49279]   :/ A_weights[769],
      [49280 : 49343]   :/ A_weights[770],
      [49344 : 49407]   :/ A_weights[771],
      [49408 : 49471]   :/ A_weights[772],
      [49472 : 49535]   :/ A_weights[773],
      [49536 : 49599]   :/ A_weights[774],
      [49600 : 49663]   :/ A_weights[775],
      [49664 : 49727]   :/ A_weights[776],
      [49728 : 49791]   :/ A_weights[777],
      [49792 : 49855]   :/ A_weights[778],
      [49856 : 49919]   :/ A_weights[779],
      [49920 : 49983]   :/ A_weights[780],
      [49984 : 50047]   :/ A_weights[781],
      [50048 : 50111]   :/ A_weights[782],
      [50112 : 50175]   :/ A_weights[783],
      [50176 : 50239]   :/ A_weights[784],
      [50240 : 50303]   :/ A_weights[785],
      [50304 : 50367]   :/ A_weights[786],
      [50368 : 50431]   :/ A_weights[787],
      [50432 : 50495]   :/ A_weights[788],
      [50496 : 50559]   :/ A_weights[789],
      [50560 : 50623]   :/ A_weights[790],
      [50624 : 50687]   :/ A_weights[791],
      [50688 : 50751]   :/ A_weights[792],
      [50752 : 50815]   :/ A_weights[793],
      [50816 : 50879]   :/ A_weights[794],
      [50880 : 50943]   :/ A_weights[795],
      [50944 : 51007]   :/ A_weights[796],
      [51008 : 51071]   :/ A_weights[797],
      [51072 : 51135]   :/ A_weights[798],
      [51136 : 51199]   :/ A_weights[799],
      [51200 : 51263]   :/ A_weights[800],
      [51264 : 51327]   :/ A_weights[801],
      [51328 : 51391]   :/ A_weights[802],
      [51392 : 51455]   :/ A_weights[803],
      [51456 : 51519]   :/ A_weights[804],
      [51520 : 51583]   :/ A_weights[805],
      [51584 : 51647]   :/ A_weights[806],
      [51648 : 51711]   :/ A_weights[807],
      [51712 : 51775]   :/ A_weights[808],
      [51776 : 51839]   :/ A_weights[809],
      [51840 : 51903]   :/ A_weights[810],
      [51904 : 51967]   :/ A_weights[811],
      [51968 : 52031]   :/ A_weights[812],
      [52032 : 52095]   :/ A_weights[813],
      [52096 : 52159]   :/ A_weights[814],
      [52160 : 52223]   :/ A_weights[815],
      [52224 : 52287]   :/ A_weights[816],
      [52288 : 52351]   :/ A_weights[817],
      [52352 : 52415]   :/ A_weights[818],
      [52416 : 52479]   :/ A_weights[819],
      [52480 : 52543]   :/ A_weights[820],
      [52544 : 52607]   :/ A_weights[821],
      [52608 : 52671]   :/ A_weights[822],
      [52672 : 52735]   :/ A_weights[823],
      [52736 : 52799]   :/ A_weights[824],
      [52800 : 52863]   :/ A_weights[825],
      [52864 : 52927]   :/ A_weights[826],
      [52928 : 52991]   :/ A_weights[827],
      [52992 : 53055]   :/ A_weights[828],
      [53056 : 53119]   :/ A_weights[829],
      [53120 : 53183]   :/ A_weights[830],
      [53184 : 53247]   :/ A_weights[831],
      [53248 : 53311]   :/ A_weights[832],
      [53312 : 53375]   :/ A_weights[833],
      [53376 : 53439]   :/ A_weights[834],
      [53440 : 53503]   :/ A_weights[835],
      [53504 : 53567]   :/ A_weights[836],
      [53568 : 53631]   :/ A_weights[837],
      [53632 : 53695]   :/ A_weights[838],
      [53696 : 53759]   :/ A_weights[839],
      [53760 : 53823]   :/ A_weights[840],
      [53824 : 53887]   :/ A_weights[841],
      [53888 : 53951]   :/ A_weights[842],
      [53952 : 54015]   :/ A_weights[843],
      [54016 : 54079]   :/ A_weights[844],
      [54080 : 54143]   :/ A_weights[845],
      [54144 : 54207]   :/ A_weights[846],
      [54208 : 54271]   :/ A_weights[847],
      [54272 : 54335]   :/ A_weights[848],
      [54336 : 54399]   :/ A_weights[849],
      [54400 : 54463]   :/ A_weights[850],
      [54464 : 54527]   :/ A_weights[851],
      [54528 : 54591]   :/ A_weights[852],
      [54592 : 54655]   :/ A_weights[853],
      [54656 : 54719]   :/ A_weights[854],
      [54720 : 54783]   :/ A_weights[855],
      [54784 : 54847]   :/ A_weights[856],
      [54848 : 54911]   :/ A_weights[857],
      [54912 : 54975]   :/ A_weights[858],
      [54976 : 55039]   :/ A_weights[859],
      [55040 : 55103]   :/ A_weights[860],
      [55104 : 55167]   :/ A_weights[861],
      [55168 : 55231]   :/ A_weights[862],
      [55232 : 55295]   :/ A_weights[863],
      [55296 : 55359]   :/ A_weights[864],
      [55360 : 55423]   :/ A_weights[865],
      [55424 : 55487]   :/ A_weights[866],
      [55488 : 55551]   :/ A_weights[867],
      [55552 : 55615]   :/ A_weights[868],
      [55616 : 55679]   :/ A_weights[869],
      [55680 : 55743]   :/ A_weights[870],
      [55744 : 55807]   :/ A_weights[871],
      [55808 : 55871]   :/ A_weights[872],
      [55872 : 55935]   :/ A_weights[873],
      [55936 : 55999]   :/ A_weights[874],
      [56000 : 56063]   :/ A_weights[875],
      [56064 : 56127]   :/ A_weights[876],
      [56128 : 56191]   :/ A_weights[877],
      [56192 : 56255]   :/ A_weights[878],
      [56256 : 56319]   :/ A_weights[879],
      [56320 : 56383]   :/ A_weights[880],
      [56384 : 56447]   :/ A_weights[881],
      [56448 : 56511]   :/ A_weights[882],
      [56512 : 56575]   :/ A_weights[883],
      [56576 : 56639]   :/ A_weights[884],
      [56640 : 56703]   :/ A_weights[885],
      [56704 : 56767]   :/ A_weights[886],
      [56768 : 56831]   :/ A_weights[887],
      [56832 : 56895]   :/ A_weights[888],
      [56896 : 56959]   :/ A_weights[889],
      [56960 : 57023]   :/ A_weights[890],
      [57024 : 57087]   :/ A_weights[891],
      [57088 : 57151]   :/ A_weights[892],
      [57152 : 57215]   :/ A_weights[893],
      [57216 : 57279]   :/ A_weights[894],
      [57280 : 57343]   :/ A_weights[895],
      [57344 : 57407]   :/ A_weights[896],
      [57408 : 57471]   :/ A_weights[897],
      [57472 : 57535]   :/ A_weights[898],
      [57536 : 57599]   :/ A_weights[899],
      [57600 : 57663]   :/ A_weights[900],
      [57664 : 57727]   :/ A_weights[901],
      [57728 : 57791]   :/ A_weights[902],
      [57792 : 57855]   :/ A_weights[903],
      [57856 : 57919]   :/ A_weights[904],
      [57920 : 57983]   :/ A_weights[905],
      [57984 : 58047]   :/ A_weights[906],
      [58048 : 58111]   :/ A_weights[907],
      [58112 : 58175]   :/ A_weights[908],
      [58176 : 58239]   :/ A_weights[909],
      [58240 : 58303]   :/ A_weights[910],
      [58304 : 58367]   :/ A_weights[911],
      [58368 : 58431]   :/ A_weights[912],
      [58432 : 58495]   :/ A_weights[913],
      [58496 : 58559]   :/ A_weights[914],
      [58560 : 58623]   :/ A_weights[915],
      [58624 : 58687]   :/ A_weights[916],
      [58688 : 58751]   :/ A_weights[917],
      [58752 : 58815]   :/ A_weights[918],
      [58816 : 58879]   :/ A_weights[919],
      [58880 : 58943]   :/ A_weights[920],
      [58944 : 59007]   :/ A_weights[921],
      [59008 : 59071]   :/ A_weights[922],
      [59072 : 59135]   :/ A_weights[923],
      [59136 : 59199]   :/ A_weights[924],
      [59200 : 59263]   :/ A_weights[925],
      [59264 : 59327]   :/ A_weights[926],
      [59328 : 59391]   :/ A_weights[927],
      [59392 : 59455]   :/ A_weights[928],
      [59456 : 59519]   :/ A_weights[929],
      [59520 : 59583]   :/ A_weights[930],
      [59584 : 59647]   :/ A_weights[931],
      [59648 : 59711]   :/ A_weights[932],
      [59712 : 59775]   :/ A_weights[933],
      [59776 : 59839]   :/ A_weights[934],
      [59840 : 59903]   :/ A_weights[935],
      [59904 : 59967]   :/ A_weights[936],
      [59968 : 60031]   :/ A_weights[937],
      [60032 : 60095]   :/ A_weights[938],
      [60096 : 60159]   :/ A_weights[939],
      [60160 : 60223]   :/ A_weights[940],
      [60224 : 60287]   :/ A_weights[941],
      [60288 : 60351]   :/ A_weights[942],
      [60352 : 60415]   :/ A_weights[943],
      [60416 : 60479]   :/ A_weights[944],
      [60480 : 60543]   :/ A_weights[945],
      [60544 : 60607]   :/ A_weights[946],
      [60608 : 60671]   :/ A_weights[947],
      [60672 : 60735]   :/ A_weights[948],
      [60736 : 60799]   :/ A_weights[949],
      [60800 : 60863]   :/ A_weights[950],
      [60864 : 60927]   :/ A_weights[951],
      [60928 : 60991]   :/ A_weights[952],
      [60992 : 61055]   :/ A_weights[953],
      [61056 : 61119]   :/ A_weights[954],
      [61120 : 61183]   :/ A_weights[955],
      [61184 : 61247]   :/ A_weights[956],
      [61248 : 61311]   :/ A_weights[957],
      [61312 : 61375]   :/ A_weights[958],
      [61376 : 61439]   :/ A_weights[959],
      [61440 : 61503]   :/ A_weights[960],
      [61504 : 61567]   :/ A_weights[961],
      [61568 : 61631]   :/ A_weights[962],
      [61632 : 61695]   :/ A_weights[963],
      [61696 : 61759]   :/ A_weights[964],
      [61760 : 61823]   :/ A_weights[965],
      [61824 : 61887]   :/ A_weights[966],
      [61888 : 61951]   :/ A_weights[967],
      [61952 : 62015]   :/ A_weights[968],
      [62016 : 62079]   :/ A_weights[969],
      [62080 : 62143]   :/ A_weights[970],
      [62144 : 62207]   :/ A_weights[971],
      [62208 : 62271]   :/ A_weights[972],
      [62272 : 62335]   :/ A_weights[973],
      [62336 : 62399]   :/ A_weights[974],
      [62400 : 62463]   :/ A_weights[975],
      [62464 : 62527]   :/ A_weights[976],
      [62528 : 62591]   :/ A_weights[977],
      [62592 : 62655]   :/ A_weights[978],
      [62656 : 62719]   :/ A_weights[979],
      [62720 : 62783]   :/ A_weights[980],
      [62784 : 62847]   :/ A_weights[981],
      [62848 : 62911]   :/ A_weights[982],
      [62912 : 62975]   :/ A_weights[983],
      [62976 : 63039]   :/ A_weights[984],
      [63040 : 63103]   :/ A_weights[985],
      [63104 : 63167]   :/ A_weights[986],
      [63168 : 63231]   :/ A_weights[987],
      [63232 : 63295]   :/ A_weights[988],
      [63296 : 63359]   :/ A_weights[989],
      [63360 : 63423]   :/ A_weights[990],
      [63424 : 63487]   :/ A_weights[991],
      [63488 : 63551]   :/ A_weights[992],
      [63552 : 63615]   :/ A_weights[993],
      [63616 : 63679]   :/ A_weights[994],
      [63680 : 63743]   :/ A_weights[995],
      [63744 : 63807]   :/ A_weights[996],
      [63808 : 63871]   :/ A_weights[997],
      [63872 : 63935]   :/ A_weights[998],
      [63936 : 63999]   :/ A_weights[999],
      [64000 : 64063]   :/ A_weights[1000],
      [64064 : 64127]   :/ A_weights[1001],
      [64128 : 64191]   :/ A_weights[1002],
      [64192 : 64255]   :/ A_weights[1003],
      [64256 : 64319]   :/ A_weights[1004],
      [64320 : 64383]   :/ A_weights[1005],
      [64384 : 64447]   :/ A_weights[1006],
      [64448 : 64511]   :/ A_weights[1007],
      [64512 : 64575]   :/ A_weights[1008],
      [64576 : 64639]   :/ A_weights[1009],
      [64640 : 64703]   :/ A_weights[1010],
      [64704 : 64767]   :/ A_weights[1011],
      [64768 : 64831]   :/ A_weights[1012],
      [64832 : 64895]   :/ A_weights[1013],
      [64896 : 64959]   :/ A_weights[1014],
      [64960 : 65023]   :/ A_weights[1015],
      [65024 : 65087]   :/ A_weights[1016],
      [65088 : 65151]   :/ A_weights[1017],
      [65152 : 65215]   :/ A_weights[1018],
      [65216 : 65279]   :/ A_weights[1019],
      [65280 : 65343]   :/ A_weights[1020],
      [65344 : 65407]   :/ A_weights[1021],
      [65408 : 65471]   :/ A_weights[1022],
      [65472 : 65535]   :/ A_weights[1023]
    };

      B dist {
      [0    : 63]       :/ B_weights[0],
      [64   : 127]      :/ B_weights[1],
      [128  : 191]      :/ B_weights[2],
      [192  : 255]      :/ B_weights[3],
      [256  : 319]      :/ B_weights[4],
      [320  : 383]      :/ B_weights[5],
      [384  : 447]      :/ B_weights[6],
      [448  : 511]      :/ B_weights[7],
      [512  : 575]      :/ B_weights[8],
      [576  : 639]      :/ B_weights[9],
      [640  : 703]      :/ B_weights[10],
      [704  : 767]      :/ B_weights[11],
      [768  : 831]      :/ B_weights[12],
      [832  : 895]      :/ B_weights[13],
      [896  : 959]      :/ B_weights[14],
      [960  : 1023]     :/ B_weights[15],
      [1024 : 1087]     :/ B_weights[16],
      [1088 : 1151]     :/ B_weights[17],
      [1152 : 1215]     :/ B_weights[18],
      [1216 : 1279]     :/ B_weights[19],
      [1280 : 1343]     :/ B_weights[20],
      [1344 : 1407]     :/ B_weights[21],
      [1408 : 1471]     :/ B_weights[22],
      [1472 : 1535]     :/ B_weights[23],
      [1536 : 1599]     :/ B_weights[24],
      [1600 : 1663]     :/ B_weights[25],
      [1664 : 1727]     :/ B_weights[26],
      [1728 : 1791]     :/ B_weights[27],
      [1792 : 1855]     :/ B_weights[28],
      [1856 : 1919]     :/ B_weights[29],
      [1920 : 1983]     :/ B_weights[30],
      [1984 : 2047]     :/ B_weights[31],
      [2048 : 2111]     :/ B_weights[32],
      [2112 : 2175]     :/ B_weights[33],
      [2176 : 2239]     :/ B_weights[34],
      [2240 : 2303]     :/ B_weights[35],
      [2304 : 2367]     :/ B_weights[36],
      [2368 : 2431]     :/ B_weights[37],
      [2432 : 2495]     :/ B_weights[38],
      [2496 : 2559]     :/ B_weights[39],
      [2560 : 2623]     :/ B_weights[40],
      [2624 : 2687]     :/ B_weights[41],
      [2688 : 2751]     :/ B_weights[42],
      [2752 : 2815]     :/ B_weights[43],
      [2816 : 2879]     :/ B_weights[44],
      [2880 : 2943]     :/ B_weights[45],
      [2944 : 3007]     :/ B_weights[46],
      [3008 : 3071]     :/ B_weights[47],
      [3072 : 3135]     :/ B_weights[48],
      [3136 : 3199]     :/ B_weights[49],
      [3200 : 3263]     :/ B_weights[50],
      [3264 : 3327]     :/ B_weights[51],
      [3328 : 3391]     :/ B_weights[52],
      [3392 : 3455]     :/ B_weights[53],
      [3456 : 3519]     :/ B_weights[54],
      [3520 : 3583]     :/ B_weights[55],
      [3584 : 3647]     :/ B_weights[56],
      [3648 : 3711]     :/ B_weights[57],
      [3712 : 3775]     :/ B_weights[58],
      [3776 : 3839]     :/ B_weights[59],
      [3840 : 3903]     :/ B_weights[60],
      [3904 : 3967]     :/ B_weights[61],
      [3968 : 4031]     :/ B_weights[62],
      [4032 : 4095]     :/ B_weights[63],
      [4096 : 4159]     :/ B_weights[64],
      [4160 : 4223]     :/ B_weights[65],
      [4224 : 4287]     :/ B_weights[66],
      [4288 : 4351]     :/ B_weights[67],
      [4352 : 4415]     :/ B_weights[68],
      [4416 : 4479]     :/ B_weights[69],
      [4480 : 4543]     :/ B_weights[70],
      [4544 : 4607]     :/ B_weights[71],
      [4608 : 4671]     :/ B_weights[72],
      [4672 : 4735]     :/ B_weights[73],
      [4736 : 4799]     :/ B_weights[74],
      [4800 : 4863]     :/ B_weights[75],
      [4864 : 4927]     :/ B_weights[76],
      [4928 : 4991]     :/ B_weights[77],
      [4992 : 5055]     :/ B_weights[78],
      [5056 : 5119]     :/ B_weights[79],
      [5120 : 5183]     :/ B_weights[80],
      [5184 : 5247]     :/ B_weights[81],
      [5248 : 5311]     :/ B_weights[82],
      [5312 : 5375]     :/ B_weights[83],
      [5376 : 5439]     :/ B_weights[84],
      [5440 : 5503]     :/ B_weights[85],
      [5504 : 5567]     :/ B_weights[86],
      [5568 : 5631]     :/ B_weights[87],
      [5632 : 5695]     :/ B_weights[88],
      [5696 : 5759]     :/ B_weights[89],
      [5760 : 5823]     :/ B_weights[90],
      [5824 : 5887]     :/ B_weights[91],
      [5888 : 5951]     :/ B_weights[92],
      [5952 : 6015]     :/ B_weights[93],
      [6016 : 6079]     :/ B_weights[94],
      [6080 : 6143]     :/ B_weights[95],
      [6144 : 6207]     :/ B_weights[96],
      [6208 : 6271]     :/ B_weights[97],
      [6272 : 6335]     :/ B_weights[98],
      [6336 : 6399]     :/ B_weights[99],
      [6400 : 6463]     :/ B_weights[100],
      [6464 : 6527]     :/ B_weights[101],
      [6528 : 6591]     :/ B_weights[102],
      [6592 : 6655]     :/ B_weights[103],
      [6656 : 6719]     :/ B_weights[104],
      [6720 : 6783]     :/ B_weights[105],
      [6784 : 6847]     :/ B_weights[106],
      [6848 : 6911]     :/ B_weights[107],
      [6912 : 6975]     :/ B_weights[108],
      [6976 : 7039]     :/ B_weights[109],
      [7040 : 7103]     :/ B_weights[110],
      [7104 : 7167]     :/ B_weights[111],
      [7168 : 7231]     :/ B_weights[112],
      [7232 : 7295]     :/ B_weights[113],
      [7296 : 7359]     :/ B_weights[114],
      [7360 : 7423]     :/ B_weights[115],
      [7424 : 7487]     :/ B_weights[116],
      [7488 : 7551]     :/ B_weights[117],
      [7552 : 7615]     :/ B_weights[118],
      [7616 : 7679]     :/ B_weights[119],
      [7680 : 7743]     :/ B_weights[120],
      [7744 : 7807]     :/ B_weights[121],
      [7808 : 7871]     :/ B_weights[122],
      [7872 : 7935]     :/ B_weights[123],
      [7936 : 7999]     :/ B_weights[124],
      [8000 : 8063]     :/ B_weights[125],
      [8064 : 8127]     :/ B_weights[126],
      [8128 : 8191]     :/ B_weights[127],
      [8192 : 8255]     :/ B_weights[128],
      [8256 : 8319]     :/ B_weights[129],
      [8320 : 8383]     :/ B_weights[130],
      [8384 : 8447]     :/ B_weights[131],
      [8448 : 8511]     :/ B_weights[132],
      [8512 : 8575]     :/ B_weights[133],
      [8576 : 8639]     :/ B_weights[134],
      [8640 : 8703]     :/ B_weights[135],
      [8704 : 8767]     :/ B_weights[136],
      [8768 : 8831]     :/ B_weights[137],
      [8832 : 8895]     :/ B_weights[138],
      [8896 : 8959]     :/ B_weights[139],
      [8960 : 9023]     :/ B_weights[140],
      [9024 : 9087]     :/ B_weights[141],
      [9088 : 9151]     :/ B_weights[142],
      [9152 : 9215]     :/ B_weights[143],
      [9216 : 9279]     :/ B_weights[144],
      [9280 : 9343]     :/ B_weights[145],
      [9344 : 9407]     :/ B_weights[146],
      [9408 : 9471]     :/ B_weights[147],
      [9472 : 9535]     :/ B_weights[148],
      [9536 : 9599]     :/ B_weights[149],
      [9600 : 9663]     :/ B_weights[150],
      [9664 : 9727]     :/ B_weights[151],
      [9728 : 9791]     :/ B_weights[152],
      [9792 : 9855]     :/ B_weights[153],
      [9856 : 9919]     :/ B_weights[154],
      [9920 : 9983]     :/ B_weights[155],
      [9984 : 10047]    :/ B_weights[156],
      [10048 : 10111]   :/ B_weights[157],
      [10112 : 10175]   :/ B_weights[158],
      [10176 : 10239]   :/ B_weights[159],
      [10240 : 10303]   :/ B_weights[160],
      [10304 : 10367]   :/ B_weights[161],
      [10368 : 10431]   :/ B_weights[162],
      [10432 : 10495]   :/ B_weights[163],
      [10496 : 10559]   :/ B_weights[164],
      [10560 : 10623]   :/ B_weights[165],
      [10624 : 10687]   :/ B_weights[166],
      [10688 : 10751]   :/ B_weights[167],
      [10752 : 10815]   :/ B_weights[168],
      [10816 : 10879]   :/ B_weights[169],
      [10880 : 10943]   :/ B_weights[170],
      [10944 : 11007]   :/ B_weights[171],
      [11008 : 11071]   :/ B_weights[172],
      [11072 : 11135]   :/ B_weights[173],
      [11136 : 11199]   :/ B_weights[174],
      [11200 : 11263]   :/ B_weights[175],
      [11264 : 11327]   :/ B_weights[176],
      [11328 : 11391]   :/ B_weights[177],
      [11392 : 11455]   :/ B_weights[178],
      [11456 : 11519]   :/ B_weights[179],
      [11520 : 11583]   :/ B_weights[180],
      [11584 : 11647]   :/ B_weights[181],
      [11648 : 11711]   :/ B_weights[182],
      [11712 : 11775]   :/ B_weights[183],
      [11776 : 11839]   :/ B_weights[184],
      [11840 : 11903]   :/ B_weights[185],
      [11904 : 11967]   :/ B_weights[186],
      [11968 : 12031]   :/ B_weights[187],
      [12032 : 12095]   :/ B_weights[188],
      [12096 : 12159]   :/ B_weights[189],
      [12160 : 12223]   :/ B_weights[190],
      [12224 : 12287]   :/ B_weights[191],
      [12288 : 12351]   :/ B_weights[192],
      [12352 : 12415]   :/ B_weights[193],
      [12416 : 12479]   :/ B_weights[194],
      [12480 : 12543]   :/ B_weights[195],
      [12544 : 12607]   :/ B_weights[196],
      [12608 : 12671]   :/ B_weights[197],
      [12672 : 12735]   :/ B_weights[198],
      [12736 : 12799]   :/ B_weights[199],
      [12800 : 12863]   :/ B_weights[200],
      [12864 : 12927]   :/ B_weights[201],
      [12928 : 12991]   :/ B_weights[202],
      [12992 : 13055]   :/ B_weights[203],
      [13056 : 13119]   :/ B_weights[204],
      [13120 : 13183]   :/ B_weights[205],
      [13184 : 13247]   :/ B_weights[206],
      [13248 : 13311]   :/ B_weights[207],
      [13312 : 13375]   :/ B_weights[208],
      [13376 : 13439]   :/ B_weights[209],
      [13440 : 13503]   :/ B_weights[210],
      [13504 : 13567]   :/ B_weights[211],
      [13568 : 13631]   :/ B_weights[212],
      [13632 : 13695]   :/ B_weights[213],
      [13696 : 13759]   :/ B_weights[214],
      [13760 : 13823]   :/ B_weights[215],
      [13824 : 13887]   :/ B_weights[216],
      [13888 : 13951]   :/ B_weights[217],
      [13952 : 14015]   :/ B_weights[218],
      [14016 : 14079]   :/ B_weights[219],
      [14080 : 14143]   :/ B_weights[220],
      [14144 : 14207]   :/ B_weights[221],
      [14208 : 14271]   :/ B_weights[222],
      [14272 : 14335]   :/ B_weights[223],
      [14336 : 14399]   :/ B_weights[224],
      [14400 : 14463]   :/ B_weights[225],
      [14464 : 14527]   :/ B_weights[226],
      [14528 : 14591]   :/ B_weights[227],
      [14592 : 14655]   :/ B_weights[228],
      [14656 : 14719]   :/ B_weights[229],
      [14720 : 14783]   :/ B_weights[230],
      [14784 : 14847]   :/ B_weights[231],
      [14848 : 14911]   :/ B_weights[232],
      [14912 : 14975]   :/ B_weights[233],
      [14976 : 15039]   :/ B_weights[234],
      [15040 : 15103]   :/ B_weights[235],
      [15104 : 15167]   :/ B_weights[236],
      [15168 : 15231]   :/ B_weights[237],
      [15232 : 15295]   :/ B_weights[238],
      [15296 : 15359]   :/ B_weights[239],
      [15360 : 15423]   :/ B_weights[240],
      [15424 : 15487]   :/ B_weights[241],
      [15488 : 15551]   :/ B_weights[242],
      [15552 : 15615]   :/ B_weights[243],
      [15616 : 15679]   :/ B_weights[244],
      [15680 : 15743]   :/ B_weights[245],
      [15744 : 15807]   :/ B_weights[246],
      [15808 : 15871]   :/ B_weights[247],
      [15872 : 15935]   :/ B_weights[248],
      [15936 : 15999]   :/ B_weights[249],
      [16000 : 16063]   :/ B_weights[250],
      [16064 : 16127]   :/ B_weights[251],
      [16128 : 16191]   :/ B_weights[252],
      [16192 : 16255]   :/ B_weights[253],
      [16256 : 16319]   :/ B_weights[254],
      [16320 : 16383]   :/ B_weights[255],
      [16384 : 16447]   :/ B_weights[256],
      [16448 : 16511]   :/ B_weights[257],
      [16512 : 16575]   :/ B_weights[258],
      [16576 : 16639]   :/ B_weights[259],
      [16640 : 16703]   :/ B_weights[260],
      [16704 : 16767]   :/ B_weights[261],
      [16768 : 16831]   :/ B_weights[262],
      [16832 : 16895]   :/ B_weights[263],
      [16896 : 16959]   :/ B_weights[264],
      [16960 : 17023]   :/ B_weights[265],
      [17024 : 17087]   :/ B_weights[266],
      [17088 : 17151]   :/ B_weights[267],
      [17152 : 17215]   :/ B_weights[268],
      [17216 : 17279]   :/ B_weights[269],
      [17280 : 17343]   :/ B_weights[270],
      [17344 : 17407]   :/ B_weights[271],
      [17408 : 17471]   :/ B_weights[272],
      [17472 : 17535]   :/ B_weights[273],
      [17536 : 17599]   :/ B_weights[274],
      [17600 : 17663]   :/ B_weights[275],
      [17664 : 17727]   :/ B_weights[276],
      [17728 : 17791]   :/ B_weights[277],
      [17792 : 17855]   :/ B_weights[278],
      [17856 : 17919]   :/ B_weights[279],
      [17920 : 17983]   :/ B_weights[280],
      [17984 : 18047]   :/ B_weights[281],
      [18048 : 18111]   :/ B_weights[282],
      [18112 : 18175]   :/ B_weights[283],
      [18176 : 18239]   :/ B_weights[284],
      [18240 : 18303]   :/ B_weights[285],
      [18304 : 18367]   :/ B_weights[286],
      [18368 : 18431]   :/ B_weights[287],
      [18432 : 18495]   :/ B_weights[288],
      [18496 : 18559]   :/ B_weights[289],
      [18560 : 18623]   :/ B_weights[290],
      [18624 : 18687]   :/ B_weights[291],
      [18688 : 18751]   :/ B_weights[292],
      [18752 : 18815]   :/ B_weights[293],
      [18816 : 18879]   :/ B_weights[294],
      [18880 : 18943]   :/ B_weights[295],
      [18944 : 19007]   :/ B_weights[296],
      [19008 : 19071]   :/ B_weights[297],
      [19072 : 19135]   :/ B_weights[298],
      [19136 : 19199]   :/ B_weights[299],
      [19200 : 19263]   :/ B_weights[300],
      [19264 : 19327]   :/ B_weights[301],
      [19328 : 19391]   :/ B_weights[302],
      [19392 : 19455]   :/ B_weights[303],
      [19456 : 19519]   :/ B_weights[304],
      [19520 : 19583]   :/ B_weights[305],
      [19584 : 19647]   :/ B_weights[306],
      [19648 : 19711]   :/ B_weights[307],
      [19712 : 19775]   :/ B_weights[308],
      [19776 : 19839]   :/ B_weights[309],
      [19840 : 19903]   :/ B_weights[310],
      [19904 : 19967]   :/ B_weights[311],
      [19968 : 20031]   :/ B_weights[312],
      [20032 : 20095]   :/ B_weights[313],
      [20096 : 20159]   :/ B_weights[314],
      [20160 : 20223]   :/ B_weights[315],
      [20224 : 20287]   :/ B_weights[316],
      [20288 : 20351]   :/ B_weights[317],
      [20352 : 20415]   :/ B_weights[318],
      [20416 : 20479]   :/ B_weights[319],
      [20480 : 20543]   :/ B_weights[320],
      [20544 : 20607]   :/ B_weights[321],
      [20608 : 20671]   :/ B_weights[322],
      [20672 : 20735]   :/ B_weights[323],
      [20736 : 20799]   :/ B_weights[324],
      [20800 : 20863]   :/ B_weights[325],
      [20864 : 20927]   :/ B_weights[326],
      [20928 : 20991]   :/ B_weights[327],
      [20992 : 21055]   :/ B_weights[328],
      [21056 : 21119]   :/ B_weights[329],
      [21120 : 21183]   :/ B_weights[330],
      [21184 : 21247]   :/ B_weights[331],
      [21248 : 21311]   :/ B_weights[332],
      [21312 : 21375]   :/ B_weights[333],
      [21376 : 21439]   :/ B_weights[334],
      [21440 : 21503]   :/ B_weights[335],
      [21504 : 21567]   :/ B_weights[336],
      [21568 : 21631]   :/ B_weights[337],
      [21632 : 21695]   :/ B_weights[338],
      [21696 : 21759]   :/ B_weights[339],
      [21760 : 21823]   :/ B_weights[340],
      [21824 : 21887]   :/ B_weights[341],
      [21888 : 21951]   :/ B_weights[342],
      [21952 : 22015]   :/ B_weights[343],
      [22016 : 22079]   :/ B_weights[344],
      [22080 : 22143]   :/ B_weights[345],
      [22144 : 22207]   :/ B_weights[346],
      [22208 : 22271]   :/ B_weights[347],
      [22272 : 22335]   :/ B_weights[348],
      [22336 : 22399]   :/ B_weights[349],
      [22400 : 22463]   :/ B_weights[350],
      [22464 : 22527]   :/ B_weights[351],
      [22528 : 22591]   :/ B_weights[352],
      [22592 : 22655]   :/ B_weights[353],
      [22656 : 22719]   :/ B_weights[354],
      [22720 : 22783]   :/ B_weights[355],
      [22784 : 22847]   :/ B_weights[356],
      [22848 : 22911]   :/ B_weights[357],
      [22912 : 22975]   :/ B_weights[358],
      [22976 : 23039]   :/ B_weights[359],
      [23040 : 23103]   :/ B_weights[360],
      [23104 : 23167]   :/ B_weights[361],
      [23168 : 23231]   :/ B_weights[362],
      [23232 : 23295]   :/ B_weights[363],
      [23296 : 23359]   :/ B_weights[364],
      [23360 : 23423]   :/ B_weights[365],
      [23424 : 23487]   :/ B_weights[366],
      [23488 : 23551]   :/ B_weights[367],
      [23552 : 23615]   :/ B_weights[368],
      [23616 : 23679]   :/ B_weights[369],
      [23680 : 23743]   :/ B_weights[370],
      [23744 : 23807]   :/ B_weights[371],
      [23808 : 23871]   :/ B_weights[372],
      [23872 : 23935]   :/ B_weights[373],
      [23936 : 23999]   :/ B_weights[374],
      [24000 : 24063]   :/ B_weights[375],
      [24064 : 24127]   :/ B_weights[376],
      [24128 : 24191]   :/ B_weights[377],
      [24192 : 24255]   :/ B_weights[378],
      [24256 : 24319]   :/ B_weights[379],
      [24320 : 24383]   :/ B_weights[380],
      [24384 : 24447]   :/ B_weights[381],
      [24448 : 24511]   :/ B_weights[382],
      [24512 : 24575]   :/ B_weights[383],
      [24576 : 24639]   :/ B_weights[384],
      [24640 : 24703]   :/ B_weights[385],
      [24704 : 24767]   :/ B_weights[386],
      [24768 : 24831]   :/ B_weights[387],
      [24832 : 24895]   :/ B_weights[388],
      [24896 : 24959]   :/ B_weights[389],
      [24960 : 25023]   :/ B_weights[390],
      [25024 : 25087]   :/ B_weights[391],
      [25088 : 25151]   :/ B_weights[392],
      [25152 : 25215]   :/ B_weights[393],
      [25216 : 25279]   :/ B_weights[394],
      [25280 : 25343]   :/ B_weights[395],
      [25344 : 25407]   :/ B_weights[396],
      [25408 : 25471]   :/ B_weights[397],
      [25472 : 25535]   :/ B_weights[398],
      [25536 : 25599]   :/ B_weights[399],
      [25600 : 25663]   :/ B_weights[400],
      [25664 : 25727]   :/ B_weights[401],
      [25728 : 25791]   :/ B_weights[402],
      [25792 : 25855]   :/ B_weights[403],
      [25856 : 25919]   :/ B_weights[404],
      [25920 : 25983]   :/ B_weights[405],
      [25984 : 26047]   :/ B_weights[406],
      [26048 : 26111]   :/ B_weights[407],
      [26112 : 26175]   :/ B_weights[408],
      [26176 : 26239]   :/ B_weights[409],
      [26240 : 26303]   :/ B_weights[410],
      [26304 : 26367]   :/ B_weights[411],
      [26368 : 26431]   :/ B_weights[412],
      [26432 : 26495]   :/ B_weights[413],
      [26496 : 26559]   :/ B_weights[414],
      [26560 : 26623]   :/ B_weights[415],
      [26624 : 26687]   :/ B_weights[416],
      [26688 : 26751]   :/ B_weights[417],
      [26752 : 26815]   :/ B_weights[418],
      [26816 : 26879]   :/ B_weights[419],
      [26880 : 26943]   :/ B_weights[420],
      [26944 : 27007]   :/ B_weights[421],
      [27008 : 27071]   :/ B_weights[422],
      [27072 : 27135]   :/ B_weights[423],
      [27136 : 27199]   :/ B_weights[424],
      [27200 : 27263]   :/ B_weights[425],
      [27264 : 27327]   :/ B_weights[426],
      [27328 : 27391]   :/ B_weights[427],
      [27392 : 27455]   :/ B_weights[428],
      [27456 : 27519]   :/ B_weights[429],
      [27520 : 27583]   :/ B_weights[430],
      [27584 : 27647]   :/ B_weights[431],
      [27648 : 27711]   :/ B_weights[432],
      [27712 : 27775]   :/ B_weights[433],
      [27776 : 27839]   :/ B_weights[434],
      [27840 : 27903]   :/ B_weights[435],
      [27904 : 27967]   :/ B_weights[436],
      [27968 : 28031]   :/ B_weights[437],
      [28032 : 28095]   :/ B_weights[438],
      [28096 : 28159]   :/ B_weights[439],
      [28160 : 28223]   :/ B_weights[440],
      [28224 : 28287]   :/ B_weights[441],
      [28288 : 28351]   :/ B_weights[442],
      [28352 : 28415]   :/ B_weights[443],
      [28416 : 28479]   :/ B_weights[444],
      [28480 : 28543]   :/ B_weights[445],
      [28544 : 28607]   :/ B_weights[446],
      [28608 : 28671]   :/ B_weights[447],
      [28672 : 28735]   :/ B_weights[448],
      [28736 : 28799]   :/ B_weights[449],
      [28800 : 28863]   :/ B_weights[450],
      [28864 : 28927]   :/ B_weights[451],
      [28928 : 28991]   :/ B_weights[452],
      [28992 : 29055]   :/ B_weights[453],
      [29056 : 29119]   :/ B_weights[454],
      [29120 : 29183]   :/ B_weights[455],
      [29184 : 29247]   :/ B_weights[456],
      [29248 : 29311]   :/ B_weights[457],
      [29312 : 29375]   :/ B_weights[458],
      [29376 : 29439]   :/ B_weights[459],
      [29440 : 29503]   :/ B_weights[460],
      [29504 : 29567]   :/ B_weights[461],
      [29568 : 29631]   :/ B_weights[462],
      [29632 : 29695]   :/ B_weights[463],
      [29696 : 29759]   :/ B_weights[464],
      [29760 : 29823]   :/ B_weights[465],
      [29824 : 29887]   :/ B_weights[466],
      [29888 : 29951]   :/ B_weights[467],
      [29952 : 30015]   :/ B_weights[468],
      [30016 : 30079]   :/ B_weights[469],
      [30080 : 30143]   :/ B_weights[470],
      [30144 : 30207]   :/ B_weights[471],
      [30208 : 30271]   :/ B_weights[472],
      [30272 : 30335]   :/ B_weights[473],
      [30336 : 30399]   :/ B_weights[474],
      [30400 : 30463]   :/ B_weights[475],
      [30464 : 30527]   :/ B_weights[476],
      [30528 : 30591]   :/ B_weights[477],
      [30592 : 30655]   :/ B_weights[478],
      [30656 : 30719]   :/ B_weights[479],
      [30720 : 30783]   :/ B_weights[480],
      [30784 : 30847]   :/ B_weights[481],
      [30848 : 30911]   :/ B_weights[482],
      [30912 : 30975]   :/ B_weights[483],
      [30976 : 31039]   :/ B_weights[484],
      [31040 : 31103]   :/ B_weights[485],
      [31104 : 31167]   :/ B_weights[486],
      [31168 : 31231]   :/ B_weights[487],
      [31232 : 31295]   :/ B_weights[488],
      [31296 : 31359]   :/ B_weights[489],
      [31360 : 31423]   :/ B_weights[490],
      [31424 : 31487]   :/ B_weights[491],
      [31488 : 31551]   :/ B_weights[492],
      [31552 : 31615]   :/ B_weights[493],
      [31616 : 31679]   :/ B_weights[494],
      [31680 : 31743]   :/ B_weights[495],
      [31744 : 31807]   :/ B_weights[496],
      [31808 : 31871]   :/ B_weights[497],
      [31872 : 31935]   :/ B_weights[498],
      [31936 : 31999]   :/ B_weights[499],
      [32000 : 32063]   :/ B_weights[500],      
      [32064 : 32127]   :/ B_weights[501],
      [32128 : 32191]   :/ B_weights[502],
      [32192 : 32255]   :/ B_weights[503],
      [32256 : 32319]   :/ B_weights[504],
      [32320 : 32383]   :/ B_weights[505],
      [32384 : 32447]   :/ B_weights[506],
      [32448 : 32511]   :/ B_weights[507],
      [32512 : 32575]   :/ B_weights[508],
      [32576 : 32639]   :/ B_weights[509],
      [32640 : 32703]   :/ B_weights[510],
      [32704 : 32767]   :/ B_weights[511],
      [32768 : 32831]   :/ B_weights[512],
      [32832 : 32895]   :/ B_weights[513],
      [32896 : 32959]   :/ B_weights[514],
      [32960 : 33023]   :/ B_weights[515],
      [33024 : 33087]   :/ B_weights[516],
      [33088 : 33151]   :/ B_weights[517],
      [33152 : 33215]   :/ B_weights[518],
      [33216 : 33279]   :/ B_weights[519],
      [33280 : 33343]   :/ B_weights[520],
      [33344 : 33407]   :/ B_weights[521],
      [33408 : 33471]   :/ B_weights[522],
      [33472 : 33535]   :/ B_weights[523],
      [33536 : 33599]   :/ B_weights[524],
      [33600 : 33663]   :/ B_weights[525],
      [33664 : 33727]   :/ B_weights[526],
      [33728 : 33791]   :/ B_weights[527],
      [33792 : 33855]   :/ B_weights[528],
      [33856 : 33919]   :/ B_weights[529],
      [33920 : 33983]   :/ B_weights[530],
      [33984 : 34047]   :/ B_weights[531],
      [34048 : 34111]   :/ B_weights[532],
      [34112 : 34175]   :/ B_weights[533],
      [34176 : 34239]   :/ B_weights[534],
      [34240 : 34303]   :/ B_weights[535],
      [34304 : 34367]   :/ B_weights[536],
      [34368 : 34431]   :/ B_weights[537],
      [34432 : 34495]   :/ B_weights[538],
      [34496 : 34559]   :/ B_weights[539],
      [34560 : 34623]   :/ B_weights[540],
      [34624 : 34687]   :/ B_weights[541],
      [34688 : 34751]   :/ B_weights[542],
      [34752 : 34815]   :/ B_weights[543],
      [34816 : 34879]   :/ B_weights[544],
      [34880 : 34943]   :/ B_weights[545],
      [34944 : 35007]   :/ B_weights[546],
      [35008 : 35071]   :/ B_weights[547],
      [35072 : 35135]   :/ B_weights[548],
      [35136 : 35199]   :/ B_weights[549],
      [35200 : 35263]   :/ B_weights[550],
      [35264 : 35327]   :/ B_weights[551],
      [35328 : 35391]   :/ B_weights[552],
      [35392 : 35455]   :/ B_weights[553],
      [35456 : 35519]   :/ B_weights[554],
      [35520 : 35583]   :/ B_weights[555],
      [35584 : 35647]   :/ B_weights[556],
      [35648 : 35711]   :/ B_weights[557],
      [35712 : 35775]   :/ B_weights[558],
      [35776 : 35839]   :/ B_weights[559],
      [35840 : 35903]   :/ B_weights[560],
      [35904 : 35967]   :/ B_weights[561],
      [35968 : 36031]   :/ B_weights[562],
      [36032 : 36095]   :/ B_weights[563],
      [36096 : 36159]   :/ B_weights[564],
      [36160 : 36223]   :/ B_weights[565],
      [36224 : 36287]   :/ B_weights[566],
      [36288 : 36351]   :/ B_weights[567],
      [36352 : 36415]   :/ B_weights[568],
      [36416 : 36479]   :/ B_weights[569],
      [36480 : 36543]   :/ B_weights[570],
      [36544 : 36607]   :/ B_weights[571],
      [36608 : 36671]   :/ B_weights[572],
      [36672 : 36735]   :/ B_weights[573],
      [36736 : 36799]   :/ B_weights[574],
      [36800 : 36863]   :/ B_weights[575],
      [36864 : 36927]   :/ B_weights[576],
      [36928 : 36991]   :/ B_weights[577],
      [36992 : 37055]   :/ B_weights[578],
      [37056 : 37119]   :/ B_weights[579],
      [37120 : 37183]   :/ B_weights[580],
      [37184 : 37247]   :/ B_weights[581],
      [37248 : 37311]   :/ B_weights[582],
      [37312 : 37375]   :/ B_weights[583],
      [37376 : 37439]   :/ B_weights[584],
      [37440 : 37503]   :/ B_weights[585],
      [37504 : 37567]   :/ B_weights[586],
      [37568 : 37631]   :/ B_weights[587],
      [37632 : 37695]   :/ B_weights[588],
      [37696 : 37759]   :/ B_weights[589],
      [37760 : 37823]   :/ B_weights[590],
      [37824 : 37887]   :/ B_weights[591],
      [37888 : 37951]   :/ B_weights[592],
      [37952 : 38015]   :/ B_weights[593],
      [38016 : 38079]   :/ B_weights[594],
      [38080 : 38143]   :/ B_weights[595],
      [38144 : 38207]   :/ B_weights[596],
      [38208 : 38271]   :/ B_weights[597],
      [38272 : 38335]   :/ B_weights[598],
      [38336 : 38399]   :/ B_weights[599],
      [38400 : 38463]   :/ B_weights[600],
      [38464 : 38527]   :/ B_weights[601],
      [38528 : 38591]   :/ B_weights[602],
      [38592 : 38655]   :/ B_weights[603],
      [38656 : 38719]   :/ B_weights[604],
      [38720 : 38783]   :/ B_weights[605],
      [38784 : 38847]   :/ B_weights[606],
      [38848 : 38911]   :/ B_weights[607],
      [38912 : 38975]   :/ B_weights[608],
      [38976 : 39039]   :/ B_weights[609],
      [39040 : 39103]   :/ B_weights[610],
      [39104 : 39167]   :/ B_weights[611],
      [39168 : 39231]   :/ B_weights[612],
      [39232 : 39295]   :/ B_weights[613],
      [39296 : 39359]   :/ B_weights[614],
      [39360 : 39423]   :/ B_weights[615],
      [39424 : 39487]   :/ B_weights[616],
      [39488 : 39551]   :/ B_weights[617],
      [39552 : 39615]   :/ B_weights[618],
      [39616 : 39679]   :/ B_weights[619],
      [39680 : 39743]   :/ B_weights[620],
      [39744 : 39807]   :/ B_weights[621],
      [39808 : 39871]   :/ B_weights[622],
      [39872 : 39935]   :/ B_weights[623],
      [39936 : 39999]   :/ B_weights[624],
      [40000 : 40063]   :/ B_weights[625],
      [40064 : 40127]   :/ B_weights[626],
      [40128 : 40191]   :/ B_weights[627],
      [40192 : 40255]   :/ B_weights[628],
      [40256 : 40319]   :/ B_weights[629],
      [40320 : 40383]   :/ B_weights[630],
      [40384 : 40447]   :/ B_weights[631],
      [40448 : 40511]   :/ B_weights[632],
      [40512 : 40575]   :/ B_weights[633],
      [40576 : 40639]   :/ B_weights[634],
      [40640 : 40703]   :/ B_weights[635],
      [40704 : 40767]   :/ B_weights[636],
      [40768 : 40831]   :/ B_weights[637],
      [40832 : 40895]   :/ B_weights[638],
      [40896 : 40959]   :/ B_weights[639],
      [40960 : 41023]   :/ B_weights[640],
      [41024 : 41087]   :/ B_weights[641],
      [41088 : 41151]   :/ B_weights[642],
      [41152 : 41215]   :/ B_weights[643],
      [41216 : 41279]   :/ B_weights[644],
      [41280 : 41343]   :/ B_weights[645],
      [41344 : 41407]   :/ B_weights[646],
      [41408 : 41471]   :/ B_weights[647],
      [41472 : 41535]   :/ B_weights[648],
      [41536 : 41599]   :/ B_weights[649],
      [41600 : 41663]   :/ B_weights[650],
      [41664 : 41727]   :/ B_weights[651],
      [41728 : 41791]   :/ B_weights[652],
      [41792 : 41855]   :/ B_weights[653],
      [41856 : 41919]   :/ B_weights[654],
      [41920 : 41983]   :/ B_weights[655],
      [41984 : 42047]   :/ B_weights[656],
      [42048 : 42111]   :/ B_weights[657],
      [42112 : 42175]   :/ B_weights[658],
      [42176 : 42239]   :/ B_weights[659],
      [42240 : 42303]   :/ B_weights[660],
      [42304 : 42367]   :/ B_weights[661],
      [42368 : 42431]   :/ B_weights[662],
      [42432 : 42495]   :/ B_weights[663],
      [42496 : 42559]   :/ B_weights[664],
      [42560 : 42623]   :/ B_weights[665],
      [42624 : 42687]   :/ B_weights[666],
      [42688 : 42751]   :/ B_weights[667],
      [42752 : 42815]   :/ B_weights[668],
      [42816 : 42879]   :/ B_weights[669],
      [42880 : 42943]   :/ B_weights[670],
      [42944 : 43007]   :/ B_weights[671],
      [43008 : 43071]   :/ B_weights[672],
      [43072 : 43135]   :/ B_weights[673],
      [43136 : 43199]   :/ B_weights[674],
      [43200 : 43263]   :/ B_weights[675],
      [43264 : 43327]   :/ B_weights[676],
      [43328 : 43391]   :/ B_weights[677],
      [43392 : 43455]   :/ B_weights[678],
      [43456 : 43519]   :/ B_weights[679],
      [43520 : 43583]   :/ B_weights[680],
      [43584 : 43647]   :/ B_weights[681],
      [43648 : 43711]   :/ B_weights[682],
      [43712 : 43775]   :/ B_weights[683],
      [43776 : 43839]   :/ B_weights[684],
      [43840 : 43903]   :/ B_weights[685],
      [43904 : 43967]   :/ B_weights[686],
      [43968 : 44031]   :/ B_weights[687],
      [44032 : 44095]   :/ B_weights[688],
      [44096 : 44159]   :/ B_weights[689],
      [44160 : 44223]   :/ B_weights[690],
      [44224 : 44287]   :/ B_weights[691],
      [44288 : 44351]   :/ B_weights[692],
      [44352 : 44415]   :/ B_weights[693],
      [44416 : 44479]   :/ B_weights[694],
      [44480 : 44543]   :/ B_weights[695],
      [44544 : 44607]   :/ B_weights[696],
      [44608 : 44671]   :/ B_weights[697],
      [44672 : 44735]   :/ B_weights[698],
      [44736 : 44799]   :/ B_weights[699],
      [44800 : 44863]   :/ B_weights[700],
      [44864 : 44927]   :/ B_weights[701],
      [44928 : 44991]   :/ B_weights[702],
      [44992 : 45055]   :/ B_weights[703],
      [45056 : 45119]   :/ B_weights[704],
      [45120 : 45183]   :/ B_weights[705],
      [45184 : 45247]   :/ B_weights[706],
      [45248 : 45311]   :/ B_weights[707],
      [45312 : 45375]   :/ B_weights[708],
      [45376 : 45439]   :/ B_weights[709],
      [45440 : 45503]   :/ B_weights[710],
      [45504 : 45567]   :/ B_weights[711],
      [45568 : 45631]   :/ B_weights[712],
      [45632 : 45695]   :/ B_weights[713],
      [45696 : 45759]   :/ B_weights[714],
      [45760 : 45823]   :/ B_weights[715],
      [45824 : 45887]   :/ B_weights[716],
      [45888 : 45951]   :/ B_weights[717],
      [45952 : 46015]   :/ B_weights[718],
      [46016 : 46079]   :/ B_weights[719],
      [46080 : 46143]   :/ B_weights[720],
      [46144 : 46207]   :/ B_weights[721],
      [46208 : 46271]   :/ B_weights[722],
      [46272 : 46335]   :/ B_weights[723],
      [46336 : 46399]   :/ B_weights[724],
      [46400 : 46463]   :/ B_weights[725],
      [46464 : 46527]   :/ B_weights[726],
      [46528 : 46591]   :/ B_weights[727],
      [46592 : 46655]   :/ B_weights[728],
      [46656 : 46719]   :/ B_weights[729],
      [46720 : 46783]   :/ B_weights[730],
      [46784 : 46847]   :/ B_weights[731],
      [46848 : 46911]   :/ B_weights[732],
      [46912 : 46975]   :/ B_weights[733],
      [46976 : 47039]   :/ B_weights[734],
      [47040 : 47103]   :/ B_weights[735],
      [47104 : 47167]   :/ B_weights[736],
      [47168 : 47231]   :/ B_weights[737],
      [47232 : 47295]   :/ B_weights[738],
      [47296 : 47359]   :/ B_weights[739],
      [47360 : 47423]   :/ B_weights[740],
      [47424 : 47487]   :/ B_weights[741],
      [47488 : 47551]   :/ B_weights[742],
      [47552 : 47615]   :/ B_weights[743],
      [47616 : 47679]   :/ B_weights[744],
      [47680 : 47743]   :/ B_weights[745],
      [47744 : 47807]   :/ B_weights[746],
      [47808 : 47871]   :/ B_weights[747],
      [47872 : 47935]   :/ B_weights[748],
      [47936 : 47999]   :/ B_weights[749],
      [48000 : 48063]   :/ B_weights[750],
      [48064 : 48127]   :/ B_weights[751],
      [48128 : 48191]   :/ B_weights[752],
      [48192 : 48255]   :/ B_weights[753],
      [48256 : 48319]   :/ B_weights[754],
      [48320 : 48383]   :/ B_weights[755],
      [48384 : 48447]   :/ B_weights[756],
      [48448 : 48511]   :/ B_weights[757],
      [48512 : 48575]   :/ B_weights[758],
      [48576 : 48639]   :/ B_weights[759],
      [48640 : 48703]   :/ B_weights[760],
      [48704 : 48767]   :/ B_weights[761],
      [48768 : 48831]   :/ B_weights[762],
      [48832 : 48895]   :/ B_weights[763],
      [48896 : 48959]   :/ B_weights[764],
      [48960 : 49023]   :/ B_weights[765],
      [49024 : 49087]   :/ B_weights[766],
      [49088 : 49151]   :/ B_weights[767],
      [49152 : 49215]   :/ B_weights[768],
      [49216 : 49279]   :/ B_weights[769],
      [49280 : 49343]   :/ B_weights[770],
      [49344 : 49407]   :/ B_weights[771],
      [49408 : 49471]   :/ B_weights[772],
      [49472 : 49535]   :/ B_weights[773],
      [49536 : 49599]   :/ B_weights[774],
      [49600 : 49663]   :/ B_weights[775],
      [49664 : 49727]   :/ B_weights[776],
      [49728 : 49791]   :/ B_weights[777],
      [49792 : 49855]   :/ B_weights[778],
      [49856 : 49919]   :/ B_weights[779],
      [49920 : 49983]   :/ B_weights[780],
      [49984 : 50047]   :/ B_weights[781],
      [50048 : 50111]   :/ B_weights[782],
      [50112 : 50175]   :/ B_weights[783],
      [50176 : 50239]   :/ B_weights[784],
      [50240 : 50303]   :/ B_weights[785],
      [50304 : 50367]   :/ B_weights[786],
      [50368 : 50431]   :/ B_weights[787],
      [50432 : 50495]   :/ B_weights[788],
      [50496 : 50559]   :/ B_weights[789],
      [50560 : 50623]   :/ B_weights[790],
      [50624 : 50687]   :/ B_weights[791],
      [50688 : 50751]   :/ B_weights[792],
      [50752 : 50815]   :/ B_weights[793],
      [50816 : 50879]   :/ B_weights[794],
      [50880 : 50943]   :/ B_weights[795],
      [50944 : 51007]   :/ B_weights[796],
      [51008 : 51071]   :/ B_weights[797],
      [51072 : 51135]   :/ B_weights[798],
      [51136 : 51199]   :/ B_weights[799],
      [51200 : 51263]   :/ B_weights[800],
      [51264 : 51327]   :/ B_weights[801],
      [51328 : 51391]   :/ B_weights[802],
      [51392 : 51455]   :/ B_weights[803],
      [51456 : 51519]   :/ B_weights[804],
      [51520 : 51583]   :/ B_weights[805],
      [51584 : 51647]   :/ B_weights[806],
      [51648 : 51711]   :/ B_weights[807],
      [51712 : 51775]   :/ B_weights[808],
      [51776 : 51839]   :/ B_weights[809],
      [51840 : 51903]   :/ B_weights[810],
      [51904 : 51967]   :/ B_weights[811],
      [51968 : 52031]   :/ B_weights[812],
      [52032 : 52095]   :/ B_weights[813],
      [52096 : 52159]   :/ B_weights[814],
      [52160 : 52223]   :/ B_weights[815],
      [52224 : 52287]   :/ B_weights[816],
      [52288 : 52351]   :/ B_weights[817],
      [52352 : 52415]   :/ B_weights[818],
      [52416 : 52479]   :/ B_weights[819],
      [52480 : 52543]   :/ B_weights[820],
      [52544 : 52607]   :/ B_weights[821],
      [52608 : 52671]   :/ B_weights[822],
      [52672 : 52735]   :/ B_weights[823],
      [52736 : 52799]   :/ B_weights[824],
      [52800 : 52863]   :/ B_weights[825],
      [52864 : 52927]   :/ B_weights[826],
      [52928 : 52991]   :/ B_weights[827],
      [52992 : 53055]   :/ B_weights[828],
      [53056 : 53119]   :/ B_weights[829],
      [53120 : 53183]   :/ B_weights[830],
      [53184 : 53247]   :/ B_weights[831],
      [53248 : 53311]   :/ B_weights[832],
      [53312 : 53375]   :/ B_weights[833],
      [53376 : 53439]   :/ B_weights[834],
      [53440 : 53503]   :/ B_weights[835],
      [53504 : 53567]   :/ B_weights[836],
      [53568 : 53631]   :/ B_weights[837],
      [53632 : 53695]   :/ B_weights[838],
      [53696 : 53759]   :/ B_weights[839],
      [53760 : 53823]   :/ B_weights[840],
      [53824 : 53887]   :/ B_weights[841],
      [53888 : 53951]   :/ B_weights[842],
      [53952 : 54015]   :/ B_weights[843],
      [54016 : 54079]   :/ B_weights[844],
      [54080 : 54143]   :/ B_weights[845],
      [54144 : 54207]   :/ B_weights[846],
      [54208 : 54271]   :/ B_weights[847],
      [54272 : 54335]   :/ B_weights[848],
      [54336 : 54399]   :/ B_weights[849],
      [54400 : 54463]   :/ B_weights[850],
      [54464 : 54527]   :/ B_weights[851],
      [54528 : 54591]   :/ B_weights[852],
      [54592 : 54655]   :/ B_weights[853],
      [54656 : 54719]   :/ B_weights[854],
      [54720 : 54783]   :/ B_weights[855],
      [54784 : 54847]   :/ B_weights[856],
      [54848 : 54911]   :/ B_weights[857],
      [54912 : 54975]   :/ B_weights[858],
      [54976 : 55039]   :/ B_weights[859],
      [55040 : 55103]   :/ B_weights[860],
      [55104 : 55167]   :/ B_weights[861],
      [55168 : 55231]   :/ B_weights[862],
      [55232 : 55295]   :/ B_weights[863],
      [55296 : 55359]   :/ B_weights[864],
      [55360 : 55423]   :/ B_weights[865],
      [55424 : 55487]   :/ B_weights[866],
      [55488 : 55551]   :/ B_weights[867],
      [55552 : 55615]   :/ B_weights[868],
      [55616 : 55679]   :/ B_weights[869],
      [55680 : 55743]   :/ B_weights[870],
      [55744 : 55807]   :/ B_weights[871],
      [55808 : 55871]   :/ B_weights[872],
      [55872 : 55935]   :/ B_weights[873],
      [55936 : 55999]   :/ B_weights[874],
      [56000 : 56063]   :/ B_weights[875],
      [56064 : 56127]   :/ B_weights[876],
      [56128 : 56191]   :/ B_weights[877],
      [56192 : 56255]   :/ B_weights[878],
      [56256 : 56319]   :/ B_weights[879],
      [56320 : 56383]   :/ B_weights[880],
      [56384 : 56447]   :/ B_weights[881],
      [56448 : 56511]   :/ B_weights[882],
      [56512 : 56575]   :/ B_weights[883],
      [56576 : 56639]   :/ B_weights[884],
      [56640 : 56703]   :/ B_weights[885],
      [56704 : 56767]   :/ B_weights[886],
      [56768 : 56831]   :/ B_weights[887],
      [56832 : 56895]   :/ B_weights[888],
      [56896 : 56959]   :/ B_weights[889],
      [56960 : 57023]   :/ B_weights[890],
      [57024 : 57087]   :/ B_weights[891],
      [57088 : 57151]   :/ B_weights[892],
      [57152 : 57215]   :/ B_weights[893],
      [57216 : 57279]   :/ B_weights[894],
      [57280 : 57343]   :/ B_weights[895],
      [57344 : 57407]   :/ B_weights[896],
      [57408 : 57471]   :/ B_weights[897],
      [57472 : 57535]   :/ B_weights[898],
      [57536 : 57599]   :/ B_weights[899],
      [57600 : 57663]   :/ B_weights[900],
      [57664 : 57727]   :/ B_weights[901],
      [57728 : 57791]   :/ B_weights[902],
      [57792 : 57855]   :/ B_weights[903],
      [57856 : 57919]   :/ B_weights[904],
      [57920 : 57983]   :/ B_weights[905],
      [57984 : 58047]   :/ B_weights[906],
      [58048 : 58111]   :/ B_weights[907],
      [58112 : 58175]   :/ B_weights[908],
      [58176 : 58239]   :/ B_weights[909],
      [58240 : 58303]   :/ B_weights[910],
      [58304 : 58367]   :/ B_weights[911],
      [58368 : 58431]   :/ B_weights[912],
      [58432 : 58495]   :/ B_weights[913],
      [58496 : 58559]   :/ B_weights[914],
      [58560 : 58623]   :/ B_weights[915],
      [58624 : 58687]   :/ B_weights[916],
      [58688 : 58751]   :/ B_weights[917],
      [58752 : 58815]   :/ B_weights[918],
      [58816 : 58879]   :/ B_weights[919],
      [58880 : 58943]   :/ B_weights[920],
      [58944 : 59007]   :/ B_weights[921],
      [59008 : 59071]   :/ B_weights[922],
      [59072 : 59135]   :/ B_weights[923],
      [59136 : 59199]   :/ B_weights[924],
      [59200 : 59263]   :/ B_weights[925],
      [59264 : 59327]   :/ B_weights[926],
      [59328 : 59391]   :/ B_weights[927],
      [59392 : 59455]   :/ B_weights[928],
      [59456 : 59519]   :/ B_weights[929],
      [59520 : 59583]   :/ B_weights[930],
      [59584 : 59647]   :/ B_weights[931],
      [59648 : 59711]   :/ B_weights[932],
      [59712 : 59775]   :/ B_weights[933],
      [59776 : 59839]   :/ B_weights[934],
      [59840 : 59903]   :/ B_weights[935],
      [59904 : 59967]   :/ B_weights[936],
      [59968 : 60031]   :/ B_weights[937],
      [60032 : 60095]   :/ B_weights[938],
      [60096 : 60159]   :/ B_weights[939],
      [60160 : 60223]   :/ B_weights[940],
      [60224 : 60287]   :/ B_weights[941],
      [60288 : 60351]   :/ B_weights[942],
      [60352 : 60415]   :/ B_weights[943],
      [60416 : 60479]   :/ B_weights[944],
      [60480 : 60543]   :/ B_weights[945],
      [60544 : 60607]   :/ B_weights[946],
      [60608 : 60671]   :/ B_weights[947],
      [60672 : 60735]   :/ B_weights[948],
      [60736 : 60799]   :/ B_weights[949],
      [60800 : 60863]   :/ B_weights[950],
      [60864 : 60927]   :/ B_weights[951],
      [60928 : 60991]   :/ B_weights[952],
      [60992 : 61055]   :/ B_weights[953],
      [61056 : 61119]   :/ B_weights[954],
      [61120 : 61183]   :/ B_weights[955],
      [61184 : 61247]   :/ B_weights[956],
      [61248 : 61311]   :/ B_weights[957],
      [61312 : 61375]   :/ B_weights[958],
      [61376 : 61439]   :/ B_weights[959],
      [61440 : 61503]   :/ B_weights[960],
      [61504 : 61567]   :/ B_weights[961],
      [61568 : 61631]   :/ B_weights[962],
      [61632 : 61695]   :/ B_weights[963],
      [61696 : 61759]   :/ B_weights[964],
      [61760 : 61823]   :/ B_weights[965],
      [61824 : 61887]   :/ B_weights[966],
      [61888 : 61951]   :/ B_weights[967],
      [61952 : 62015]   :/ B_weights[968],
      [62016 : 62079]   :/ B_weights[969],
      [62080 : 62143]   :/ B_weights[970],
      [62144 : 62207]   :/ B_weights[971],
      [62208 : 62271]   :/ B_weights[972],
      [62272 : 62335]   :/ B_weights[973],
      [62336 : 62399]   :/ B_weights[974],
      [62400 : 62463]   :/ B_weights[975],
      [62464 : 62527]   :/ B_weights[976],
      [62528 : 62591]   :/ B_weights[977],
      [62592 : 62655]   :/ B_weights[978],
      [62656 : 62719]   :/ B_weights[979],
      [62720 : 62783]   :/ B_weights[980],
      [62784 : 62847]   :/ B_weights[981],
      [62848 : 62911]   :/ B_weights[982],
      [62912 : 62975]   :/ B_weights[983],
      [62976 : 63039]   :/ B_weights[984],
      [63040 : 63103]   :/ B_weights[985],
      [63104 : 63167]   :/ B_weights[986],
      [63168 : 63231]   :/ B_weights[987],
      [63232 : 63295]   :/ B_weights[988],
      [63296 : 63359]   :/ B_weights[989],
      [63360 : 63423]   :/ B_weights[990],
      [63424 : 63487]   :/ B_weights[991],
      [63488 : 63551]   :/ B_weights[992],
      [63552 : 63615]   :/ B_weights[993],
      [63616 : 63679]   :/ B_weights[994],
      [63680 : 63743]   :/ B_weights[995],
      [63744 : 63807]   :/ B_weights[996],
      [63808 : 63871]   :/ B_weights[997],
      [63872 : 63935]   :/ B_weights[998],
      [63936 : 63999]   :/ B_weights[999],
      [64000 : 64063]   :/ B_weights[1000],
      [64064 : 64127]   :/ B_weights[1001],
      [64128 : 64191]   :/ B_weights[1002],
      [64192 : 64255]   :/ B_weights[1003],
      [64256 : 64319]   :/ B_weights[1004],
      [64320 : 64383]   :/ B_weights[1005],
      [64384 : 64447]   :/ B_weights[1006],
      [64448 : 64511]   :/ B_weights[1007],
      [64512 : 64575]   :/ B_weights[1008],
      [64576 : 64639]   :/ B_weights[1009],
      [64640 : 64703]   :/ B_weights[1010],
      [64704 : 64767]   :/ B_weights[1011],
      [64768 : 64831]   :/ B_weights[1012],
      [64832 : 64895]   :/ B_weights[1013],
      [64896 : 64959]   :/ B_weights[1014],
      [64960 : 65023]   :/ B_weights[1015],
      [65024 : 65087]   :/ B_weights[1016],
      [65088 : 65151]   :/ B_weights[1017],
      [65152 : 65215]   :/ B_weights[1018],
      [65216 : 65279]   :/ B_weights[1019],
      [65280 : 65343]   :/ B_weights[1020],
      [65344 : 65407]   :/ B_weights[1021],
      [65408 : 65471]   :/ B_weights[1022],
      [65472 : 65535]   :/ B_weights[1023]
    };

}


