`define N 16
`define bin_count 1024
`define DEFAULT_WEIGHT 100
`define penalty 100
`define test_case_count 750